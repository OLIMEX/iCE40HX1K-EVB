// ******************************************************************************

// iCEcube Netlister

// Version:            2015.08.27744

// Build Date:         Oct 14 2015 00:55:30

// File Generated:     Jul 18 2016 09:41:18

// Purpose:            Post-Route Verilog/VHDL netlist for timing simulation

// Copyright (C) 2006-2010 by Lattice Semiconductor Corp. All rights reserved.

// ******************************************************************************

// Verilog file for cell "led_but_ex1" view "INTERFACE"

module led_but_ex1 (
    LED2,
    CLK,
    BUT1,
    LED1,
    BUT2);

    output LED2;
    input CLK;
    input BUT1;
    output LED1;
    input BUT2;

    wire N__2577;
    wire N__2576;
    wire N__2575;
    wire N__2566;
    wire N__2565;
    wire N__2564;
    wire N__2557;
    wire N__2556;
    wire N__2555;
    wire N__2548;
    wire N__2547;
    wire N__2546;
    wire N__2539;
    wire N__2538;
    wire N__2537;
    wire N__2520;
    wire N__2519;
    wire N__2516;
    wire N__2513;
    wire N__2510;
    wire N__2505;
    wire N__2502;
    wire N__2501;
    wire N__2498;
    wire N__2495;
    wire N__2492;
    wire N__2487;
    wire N__2484;
    wire N__2483;
    wire N__2480;
    wire N__2477;
    wire N__2474;
    wire N__2469;
    wire N__2466;
    wire N__2465;
    wire N__2462;
    wire N__2459;
    wire N__2456;
    wire N__2451;
    wire N__2448;
    wire N__2447;
    wire N__2444;
    wire N__2441;
    wire N__2438;
    wire N__2433;
    wire N__2430;
    wire N__2427;
    wire N__2426;
    wire N__2423;
    wire N__2420;
    wire N__2415;
    wire N__2412;
    wire N__2409;
    wire N__2406;
    wire N__2403;
    wire N__2400;
    wire N__2397;
    wire N__2396;
    wire N__2393;
    wire N__2390;
    wire N__2387;
    wire N__2382;
    wire N__2381;
    wire N__2380;
    wire N__2379;
    wire N__2378;
    wire N__2377;
    wire N__2376;
    wire N__2375;
    wire N__2374;
    wire N__2373;
    wire N__2372;
    wire N__2371;
    wire N__2370;
    wire N__2369;
    wire N__2368;
    wire N__2337;
    wire N__2334;
    wire N__2331;
    wire N__2330;
    wire N__2329;
    wire N__2328;
    wire N__2327;
    wire N__2326;
    wire N__2325;
    wire N__2324;
    wire N__2323;
    wire N__2322;
    wire N__2321;
    wire N__2320;
    wire N__2319;
    wire N__2318;
    wire N__2317;
    wire N__2316;
    wire N__2315;
    wire N__2314;
    wire N__2305;
    wire N__2298;
    wire N__2289;
    wire N__2282;
    wire N__2277;
    wire N__2272;
    wire N__2271;
    wire N__2270;
    wire N__2269;
    wire N__2268;
    wire N__2267;
    wire N__2266;
    wire N__2263;
    wire N__2260;
    wire N__2257;
    wire N__2254;
    wire N__2251;
    wire N__2248;
    wire N__2223;
    wire N__2220;
    wire N__2217;
    wire N__2214;
    wire N__2211;
    wire N__2210;
    wire N__2207;
    wire N__2204;
    wire N__2201;
    wire N__2196;
    wire N__2193;
    wire N__2192;
    wire N__2189;
    wire N__2186;
    wire N__2181;
    wire N__2178;
    wire N__2175;
    wire N__2172;
    wire N__2169;
    wire N__2166;
    wire N__2163;
    wire N__2160;
    wire N__2157;
    wire N__2154;
    wire N__2151;
    wire N__2148;
    wire N__2147;
    wire N__2144;
    wire N__2141;
    wire N__2138;
    wire N__2133;
    wire N__2132;
    wire N__2131;
    wire N__2128;
    wire N__2125;
    wire N__2122;
    wire N__2115;
    wire N__2114;
    wire N__2113;
    wire N__2112;
    wire N__2109;
    wire N__2106;
    wire N__2101;
    wire N__2098;
    wire N__2095;
    wire N__2088;
    wire N__2087;
    wire N__2084;
    wire N__2081;
    wire N__2078;
    wire N__2073;
    wire N__2070;
    wire N__2069;
    wire N__2066;
    wire N__2063;
    wire N__2060;
    wire N__2055;
    wire N__2052;
    wire N__2051;
    wire N__2048;
    wire N__2045;
    wire N__2042;
    wire N__2037;
    wire N__2034;
    wire N__2031;
    wire N__2028;
    wire N__2025;
    wire N__2024;
    wire N__2021;
    wire N__2018;
    wire N__2013;
    wire N__2010;
    wire N__2009;
    wire N__2008;
    wire N__2005;
    wire N__2000;
    wire N__1995;
    wire N__1992;
    wire N__1989;
    wire N__1986;
    wire N__1983;
    wire N__1982;
    wire N__1981;
    wire N__1980;
    wire N__1977;
    wire N__1974;
    wire N__1971;
    wire N__1968;
    wire N__1959;
    wire N__1956;
    wire N__1955;
    wire N__1952;
    wire N__1949;
    wire N__1944;
    wire N__1941;
    wire N__1938;
    wire N__1935;
    wire N__1932;
    wire N__1929;
    wire N__1928;
    wire N__1923;
    wire N__1920;
    wire N__1917;
    wire N__1916;
    wire N__1913;
    wire N__1910;
    wire N__1905;
    wire N__1902;
    wire N__1901;
    wire N__1898;
    wire N__1895;
    wire N__1890;
    wire N__1887;
    wire N__1884;
    wire N__1881;
    wire N__1878;
    wire N__1875;
    wire N__1872;
    wire N__1869;
    wire N__1866;
    wire N__1863;
    wire N__1860;
    wire N__1857;
    wire N__1854;
    wire N__1851;
    wire N__1848;
    wire N__1845;
    wire N__1842;
    wire N__1839;
    wire N__1836;
    wire N__1833;
    wire N__1830;
    wire N__1827;
    wire N__1824;
    wire N__1821;
    wire N__1818;
    wire N__1815;
    wire N__1812;
    wire N__1809;
    wire N__1806;
    wire N__1803;
    wire N__1800;
    wire N__1797;
    wire N__1796;
    wire N__1793;
    wire N__1790;
    wire N__1789;
    wire N__1784;
    wire N__1781;
    wire N__1778;
    wire N__1773;
    wire N__1770;
    wire N__1767;
    wire N__1766;
    wire N__1765;
    wire N__1762;
    wire N__1759;
    wire N__1756;
    wire N__1749;
    wire N__1748;
    wire N__1745;
    wire N__1744;
    wire N__1743;
    wire N__1742;
    wire N__1741;
    wire N__1738;
    wire N__1737;
    wire N__1736;
    wire N__1735;
    wire N__1734;
    wire N__1733;
    wire N__1730;
    wire N__1725;
    wire N__1722;
    wire N__1719;
    wire N__1714;
    wire N__1709;
    wire N__1704;
    wire N__1697;
    wire N__1694;
    wire N__1683;
    wire N__1680;
    wire N__1677;
    wire N__1676;
    wire N__1675;
    wire N__1672;
    wire N__1671;
    wire N__1668;
    wire N__1665;
    wire N__1664;
    wire N__1663;
    wire N__1662;
    wire N__1655;
    wire N__1652;
    wire N__1649;
    wire N__1646;
    wire N__1645;
    wire N__1642;
    wire N__1641;
    wire N__1636;
    wire N__1627;
    wire N__1624;
    wire N__1621;
    wire N__1614;
    wire N__1611;
    wire N__1610;
    wire N__1609;
    wire N__1608;
    wire N__1607;
    wire N__1606;
    wire N__1605;
    wire N__1604;
    wire N__1603;
    wire N__1600;
    wire N__1593;
    wire N__1584;
    wire N__1581;
    wire N__1572;
    wire N__1571;
    wire N__1570;
    wire N__1567;
    wire N__1562;
    wire N__1557;
    wire N__1556;
    wire N__1553;
    wire N__1550;
    wire N__1547;
    wire N__1542;
    wire N__1539;
    wire N__1536;
    wire N__1533;
    wire N__1530;
    wire N__1527;
    wire N__1524;
    wire N__1521;
    wire N__1518;
    wire N__1515;
    wire N__1512;
    wire N__1509;
    wire N__1506;
    wire N__1503;
    wire N__1500;
    wire N__1497;
    wire N__1496;
    wire N__1495;
    wire N__1492;
    wire N__1487;
    wire N__1482;
    wire N__1479;
    wire N__1476;
    wire N__1473;
    wire N__1470;
    wire N__1467;
    wire N__1464;
    wire N__1461;
    wire N__1460;
    wire N__1457;
    wire N__1454;
    wire N__1451;
    wire N__1446;
    wire N__1445;
    wire N__1442;
    wire N__1439;
    wire N__1436;
    wire N__1431;
    wire N__1430;
    wire N__1427;
    wire N__1424;
    wire N__1419;
    wire N__1418;
    wire N__1417;
    wire N__1414;
    wire N__1409;
    wire N__1404;
    wire N__1403;
    wire N__1402;
    wire N__1401;
    wire N__1398;
    wire N__1395;
    wire N__1390;
    wire N__1383;
    wire N__1382;
    wire N__1379;
    wire N__1378;
    wire N__1377;
    wire N__1372;
    wire N__1369;
    wire N__1366;
    wire N__1363;
    wire N__1356;
    wire N__1355;
    wire N__1354;
    wire N__1351;
    wire N__1346;
    wire N__1341;
    wire N__1338;
    wire N__1335;
    wire N__1332;
    wire N__1329;
    wire N__1328;
    wire N__1327;
    wire N__1324;
    wire N__1319;
    wire N__1314;
    wire N__1313;
    wire N__1312;
    wire N__1311;
    wire N__1306;
    wire N__1303;
    wire N__1300;
    wire N__1293;
    wire N__1292;
    wire N__1289;
    wire N__1288;
    wire N__1285;
    wire N__1282;
    wire N__1279;
    wire N__1272;
    wire N__1269;
    wire N__1266;
    wire N__1263;
    wire N__1260;
    wire N__1257;
    wire N__1256;
    wire N__1251;
    wire N__1248;
    wire N__1245;
    wire N__1242;
    wire N__1239;
    wire N__1236;
    wire N__1233;
    wire N__1230;
    wire N__1227;
    wire N__1224;
    wire N__1221;
    wire N__1218;
    wire N__1215;
    wire N__1212;
    wire N__1209;
    wire N__1206;
    wire N__1203;
    wire N__1200;
    wire N__1197;
    wire N__1194;
    wire N__1191;
    wire N__1188;
    wire VCCG0;
    wire bfn_1_4_0_;
    wire cntr_1_cry_1;
    wire cntr_1_cry_2;
    wire cntr_1_cry_3;
    wire cntr_1_5;
    wire cntr_1_cry_4;
    wire cntr_1_6;
    wire cntr_1_cry_5;
    wire cntr_1_cry_6;
    wire cntr_1_8;
    wire cntr_1_cry_7;
    wire cntr_1_cry_8;
    wire bfn_1_5_0_;
    wire cntr_1_cry_9;
    wire cntr_1_cry_10;
    wire cntr_1_cry_11;
    wire cntr_1_cry_12;
    wire cntr_1_cry_13;
    wire clk_div_RNIM1KP1Z0Z_11;
    wire BUT1_r_RNIKV9MZ0Z2_cascade_;
    wire cntr_RNITQ4V2Z0Z_14;
    wire LED1_m1_r_cnv_7_cascade_;
    wire cntr_RNIV9NN2Z0Z_4;
    wire cntr7lto7_0_4_cascade_;
    wire cntrZ0Z_8;
    wire LED1_m1_r_cnv_5;
    wire LED1_m1_r_cnv_6;
    wire cntr7lto7_0_2;
    wire cntrZ0Z_2;
    wire cntrZ0Z_3;
    wire cntr7lt5_3;
    wire cntrZ0Z_6;
    wire cntrZ0Z_5;
    wire cntrZ0Z_7;
    wire cntrZ0Z_4;
    wire cntr7lto7_c;
    wire cntr_1_10;
    wire cntrZ0Z_10;
    wire cntrZ0Z_0;
    wire cntrZ0Z_1;
    wire cntr_1_9;
    wire cntrZ0Z_9;
    wire cntr_1_11;
    wire cntrZ0Z_11;
    wire cntrZ0Z_13;
    wire cntr_1_12;
    wire cntrZ0Z_14;
    wire cntr7lt13;
    wire cntrZ0Z_12;
    wire rst_cnt_i_14;
    wire rst_cntZ0Z_0;
    wire bfn_2_7_0_;
    wire rst_cntZ0Z_1;
    wire un1_rst_cnt_1_cry_0;
    wire rst_cntZ0Z_2;
    wire un1_rst_cnt_1_cry_1;
    wire rst_cntZ0Z_3;
    wire un1_rst_cnt_1_cry_2;
    wire rst_cntZ0Z_4;
    wire un1_rst_cnt_1_cry_3;
    wire rst_cntZ0Z_5;
    wire un1_rst_cnt_1_cry_4;
    wire rst_cntZ0Z_6;
    wire un1_rst_cnt_1_cry_5;
    wire rst_cntZ0Z_7;
    wire un1_rst_cnt_1_cry_6;
    wire un1_rst_cnt_1_cry_7;
    wire rst_cntZ0Z_8;
    wire bfn_2_8_0_;
    wire rst_cntZ0Z_9;
    wire un1_rst_cnt_1_cry_8;
    wire rst_cntZ0Z_10;
    wire un1_rst_cnt_1_cry_9;
    wire rst_cntZ0Z_11;
    wire un1_rst_cnt_1_cry_10;
    wire rst_cntZ0Z_12;
    wire un1_rst_cnt_1_cry_11;
    wire rst_cntZ0Z_13;
    wire un1_rst_cnt_1_cry_12;
    wire un1_rst_cnt_1_cry_13;
    wire CONSTANT_ONE_NET;
    wire GNDG0;
    wire un1_rst_cnt_1_cry_13_THRU_CRY_0_THRU_CO;
    wire un1_rst_cnt_1_cry_13_THRU_CRY_1_THRU_CO;
    wire bfn_2_9_0_;
    wire rst_cntZ0Z_14;
    wire N_16_0;
    wire BUT1_r_RNIKV9MZ0Z2;
    wire LED2_m1_rZ0;
    wire LED2_c;
    wire modeZ0;
    wire LED1_m1_rZ0;
    wire LED1_c;
    wire bfn_4_7_0_;
    wire clk_div_2_cry_1;
    wire clk_div_2_cry_2;
    wire clk_div_2_cry_3;
    wire clk_div_2_cry_4;
    wire clk_div_2_cry_5;
    wire clk_div_2_cry_6;
    wire clk_div_2_cry_7;
    wire clk_div_2_cry_8;
    wire bfn_4_8_0_;
    wire clk_div_2_cry_9;
    wire clk_div_2_cry_10;
    wire clk_div_RNI06L91Z0Z_11;
    wire clk_div_i_11;
    wire LED1_m0_rZ0;
    wire LED2_m0_rZ0;
    wire BUT2_c;
    wire BUT2_rZ0;
    wire clk_divZ0Z_1;
    wire clk_divZ0Z_0;
    wire bfn_5_7_0_;
    wire clk_divZ0Z_2;
    wire clk_div_1_cry_1;
    wire clk_divZ0Z_3;
    wire clk_div_1_cry_2;
    wire clk_divZ0Z_4;
    wire clk_div_1_cry_3;
    wire clk_divZ0Z_5;
    wire clk_div_1_cry_4;
    wire clk_divZ0Z_6;
    wire clk_div_1_cry_5;
    wire clk_divZ0Z_7;
    wire clk_div_1_cry_6;
    wire clk_divZ0Z_8;
    wire clk_div_1_cry_7;
    wire clk_div_1_cry_8;
    wire clk_divZ0Z_9;
    wire bfn_5_8_0_;
    wire clk_div_1_cry_9;
    wire clk_divZ0Z_10;
    wire BUT1_c;
    wire BUT1_rZ0;
    wire CLK_c_g;
    wire N_16_g;
    wire _gnd_net_;

    PRE_IO_GBUF CLK_ibuf_gb_io_preiogbuf (
            .PADSIGNALTOGLOBALBUFFER(N__2575),
            .GLOBALBUFFEROUTPUT(CLK_c_g));
    IO_PAD CLK_ibuf_gb_io_iopad (
            .OE(N__2577),
            .DIN(N__2576),
            .DOUT(N__2575),
            .PACKAGEPIN(CLK));
    defparam CLK_ibuf_gb_io_preio.NEG_TRIGGER=1'b0;
    defparam CLK_ibuf_gb_io_preio.PIN_TYPE=6'b000001;
    PRE_IO CLK_ibuf_gb_io_preio (
            .PADOEN(N__2577),
            .PADOUT(N__2576),
            .PADIN(N__2575),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUT2_ibuf_iopad (
            .OE(N__2566),
            .DIN(N__2565),
            .DOUT(N__2564),
            .PACKAGEPIN(BUT2));
    defparam BUT2_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam BUT2_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO BUT2_ibuf_preio (
            .PADOEN(N__2566),
            .PADOUT(N__2565),
            .PADIN(N__2564),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(BUT2_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD BUT1_ibuf_iopad (
            .OE(N__2557),
            .DIN(N__2556),
            .DOUT(N__2555),
            .PACKAGEPIN(BUT1));
    defparam BUT1_ibuf_preio.NEG_TRIGGER=1'b0;
    defparam BUT1_ibuf_preio.PIN_TYPE=6'b000001;
    PRE_IO BUT1_ibuf_preio (
            .PADOEN(N__2557),
            .PADOUT(N__2556),
            .PADIN(N__2555),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(BUT1_c),
            .DOUT0(),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LED1_obuf_iopad (
            .OE(N__2548),
            .DIN(N__2547),
            .DOUT(N__2546),
            .PACKAGEPIN(LED1));
    defparam LED1_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LED1_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LED1_obuf_preio (
            .PADOEN(N__2548),
            .PADOUT(N__2547),
            .PADIN(N__2546),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1890),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    IO_PAD LED2_obuf_iopad (
            .OE(N__2539),
            .DIN(N__2538),
            .DOUT(N__2537),
            .PACKAGEPIN(LED2));
    defparam LED2_obuf_preio.NEG_TRIGGER=1'b0;
    defparam LED2_obuf_preio.PIN_TYPE=6'b011001;
    PRE_IO LED2_obuf_preio (
            .PADOEN(N__2539),
            .PADOUT(N__2538),
            .PADIN(N__2537),
            .CLOCKENABLE(),
            .DOUT1(),
            .OUTPUTENABLE(),
            .DIN0(),
            .DOUT0(N__1944),
            .INPUTCLK(),
            .LATCHINPUTVALUE(),
            .DIN1(),
            .OUTPUTCLK());
    CascadeMux I__550 (
            .O(N__2520),
            .I(N__2516));
    InMux I__549 (
            .O(N__2519),
            .I(N__2513));
    InMux I__548 (
            .O(N__2516),
            .I(N__2510));
    LocalMux I__547 (
            .O(N__2513),
            .I(clk_divZ0Z_5));
    LocalMux I__546 (
            .O(N__2510),
            .I(clk_divZ0Z_5));
    InMux I__545 (
            .O(N__2505),
            .I(clk_div_1_cry_4));
    CascadeMux I__544 (
            .O(N__2502),
            .I(N__2498));
    InMux I__543 (
            .O(N__2501),
            .I(N__2495));
    InMux I__542 (
            .O(N__2498),
            .I(N__2492));
    LocalMux I__541 (
            .O(N__2495),
            .I(clk_divZ0Z_6));
    LocalMux I__540 (
            .O(N__2492),
            .I(clk_divZ0Z_6));
    InMux I__539 (
            .O(N__2487),
            .I(clk_div_1_cry_5));
    CascadeMux I__538 (
            .O(N__2484),
            .I(N__2480));
    InMux I__537 (
            .O(N__2483),
            .I(N__2477));
    InMux I__536 (
            .O(N__2480),
            .I(N__2474));
    LocalMux I__535 (
            .O(N__2477),
            .I(clk_divZ0Z_7));
    LocalMux I__534 (
            .O(N__2474),
            .I(clk_divZ0Z_7));
    InMux I__533 (
            .O(N__2469),
            .I(clk_div_1_cry_6));
    CascadeMux I__532 (
            .O(N__2466),
            .I(N__2462));
    InMux I__531 (
            .O(N__2465),
            .I(N__2459));
    InMux I__530 (
            .O(N__2462),
            .I(N__2456));
    LocalMux I__529 (
            .O(N__2459),
            .I(clk_divZ0Z_8));
    LocalMux I__528 (
            .O(N__2456),
            .I(clk_divZ0Z_8));
    InMux I__527 (
            .O(N__2451),
            .I(clk_div_1_cry_7));
    CascadeMux I__526 (
            .O(N__2448),
            .I(N__2444));
    InMux I__525 (
            .O(N__2447),
            .I(N__2441));
    InMux I__524 (
            .O(N__2444),
            .I(N__2438));
    LocalMux I__523 (
            .O(N__2441),
            .I(clk_divZ0Z_9));
    LocalMux I__522 (
            .O(N__2438),
            .I(clk_divZ0Z_9));
    InMux I__521 (
            .O(N__2433),
            .I(bfn_5_8_0_));
    InMux I__520 (
            .O(N__2430),
            .I(clk_div_1_cry_9));
    InMux I__519 (
            .O(N__2427),
            .I(N__2423));
    InMux I__518 (
            .O(N__2426),
            .I(N__2420));
    LocalMux I__517 (
            .O(N__2423),
            .I(clk_divZ0Z_10));
    LocalMux I__516 (
            .O(N__2420),
            .I(clk_divZ0Z_10));
    InMux I__515 (
            .O(N__2415),
            .I(N__2412));
    LocalMux I__514 (
            .O(N__2412),
            .I(N__2409));
    Span4Mux_h I__513 (
            .O(N__2409),
            .I(N__2406));
    Odrv4 I__512 (
            .O(N__2406),
            .I(BUT1_c));
    InMux I__511 (
            .O(N__2403),
            .I(N__2400));
    LocalMux I__510 (
            .O(N__2400),
            .I(N__2397));
    Span4Mux_v I__509 (
            .O(N__2397),
            .I(N__2393));
    InMux I__508 (
            .O(N__2396),
            .I(N__2390));
    Span4Mux_h I__507 (
            .O(N__2393),
            .I(N__2387));
    LocalMux I__506 (
            .O(N__2390),
            .I(BUT1_rZ0));
    Odrv4 I__505 (
            .O(N__2387),
            .I(BUT1_rZ0));
    ClkMux I__504 (
            .O(N__2382),
            .I(N__2337));
    ClkMux I__503 (
            .O(N__2381),
            .I(N__2337));
    ClkMux I__502 (
            .O(N__2380),
            .I(N__2337));
    ClkMux I__501 (
            .O(N__2379),
            .I(N__2337));
    ClkMux I__500 (
            .O(N__2378),
            .I(N__2337));
    ClkMux I__499 (
            .O(N__2377),
            .I(N__2337));
    ClkMux I__498 (
            .O(N__2376),
            .I(N__2337));
    ClkMux I__497 (
            .O(N__2375),
            .I(N__2337));
    ClkMux I__496 (
            .O(N__2374),
            .I(N__2337));
    ClkMux I__495 (
            .O(N__2373),
            .I(N__2337));
    ClkMux I__494 (
            .O(N__2372),
            .I(N__2337));
    ClkMux I__493 (
            .O(N__2371),
            .I(N__2337));
    ClkMux I__492 (
            .O(N__2370),
            .I(N__2337));
    ClkMux I__491 (
            .O(N__2369),
            .I(N__2337));
    ClkMux I__490 (
            .O(N__2368),
            .I(N__2337));
    GlobalMux I__489 (
            .O(N__2337),
            .I(N__2334));
    gio2CtrlBuf I__488 (
            .O(N__2334),
            .I(CLK_c_g));
    InMux I__487 (
            .O(N__2331),
            .I(N__2305));
    InMux I__486 (
            .O(N__2330),
            .I(N__2305));
    InMux I__485 (
            .O(N__2329),
            .I(N__2305));
    InMux I__484 (
            .O(N__2328),
            .I(N__2305));
    InMux I__483 (
            .O(N__2327),
            .I(N__2298));
    InMux I__482 (
            .O(N__2326),
            .I(N__2298));
    InMux I__481 (
            .O(N__2325),
            .I(N__2298));
    InMux I__480 (
            .O(N__2324),
            .I(N__2289));
    InMux I__479 (
            .O(N__2323),
            .I(N__2289));
    InMux I__478 (
            .O(N__2322),
            .I(N__2289));
    InMux I__477 (
            .O(N__2321),
            .I(N__2289));
    InMux I__476 (
            .O(N__2320),
            .I(N__2282));
    InMux I__475 (
            .O(N__2319),
            .I(N__2282));
    InMux I__474 (
            .O(N__2318),
            .I(N__2282));
    InMux I__473 (
            .O(N__2317),
            .I(N__2277));
    InMux I__472 (
            .O(N__2316),
            .I(N__2277));
    InMux I__471 (
            .O(N__2315),
            .I(N__2272));
    InMux I__470 (
            .O(N__2314),
            .I(N__2272));
    LocalMux I__469 (
            .O(N__2305),
            .I(N__2263));
    LocalMux I__468 (
            .O(N__2298),
            .I(N__2260));
    LocalMux I__467 (
            .O(N__2289),
            .I(N__2257));
    LocalMux I__466 (
            .O(N__2282),
            .I(N__2254));
    LocalMux I__465 (
            .O(N__2277),
            .I(N__2251));
    LocalMux I__464 (
            .O(N__2272),
            .I(N__2248));
    CEMux I__463 (
            .O(N__2271),
            .I(N__2223));
    CEMux I__462 (
            .O(N__2270),
            .I(N__2223));
    CEMux I__461 (
            .O(N__2269),
            .I(N__2223));
    CEMux I__460 (
            .O(N__2268),
            .I(N__2223));
    CEMux I__459 (
            .O(N__2267),
            .I(N__2223));
    CEMux I__458 (
            .O(N__2266),
            .I(N__2223));
    Glb2LocalMux I__457 (
            .O(N__2263),
            .I(N__2223));
    Glb2LocalMux I__456 (
            .O(N__2260),
            .I(N__2223));
    Glb2LocalMux I__455 (
            .O(N__2257),
            .I(N__2223));
    Glb2LocalMux I__454 (
            .O(N__2254),
            .I(N__2223));
    Glb2LocalMux I__453 (
            .O(N__2251),
            .I(N__2223));
    Glb2LocalMux I__452 (
            .O(N__2248),
            .I(N__2223));
    GlobalMux I__451 (
            .O(N__2223),
            .I(N__2220));
    gio2CtrlBuf I__450 (
            .O(N__2220),
            .I(N_16_g));
    InMux I__449 (
            .O(N__2217),
            .I(clk_div_2_cry_10));
    CascadeMux I__448 (
            .O(N__2214),
            .I(N__2211));
    InMux I__447 (
            .O(N__2211),
            .I(N__2207));
    InMux I__446 (
            .O(N__2210),
            .I(N__2204));
    LocalMux I__445 (
            .O(N__2207),
            .I(N__2201));
    LocalMux I__444 (
            .O(N__2204),
            .I(clk_div_RNI06L91Z0Z_11));
    Odrv4 I__443 (
            .O(N__2201),
            .I(clk_div_RNI06L91Z0Z_11));
    InMux I__442 (
            .O(N__2196),
            .I(N__2193));
    LocalMux I__441 (
            .O(N__2193),
            .I(N__2189));
    InMux I__440 (
            .O(N__2192),
            .I(N__2186));
    Odrv4 I__439 (
            .O(N__2189),
            .I(clk_div_i_11));
    LocalMux I__438 (
            .O(N__2186),
            .I(clk_div_i_11));
    InMux I__437 (
            .O(N__2181),
            .I(N__2178));
    LocalMux I__436 (
            .O(N__2178),
            .I(LED1_m0_rZ0));
    InMux I__435 (
            .O(N__2175),
            .I(N__2172));
    LocalMux I__434 (
            .O(N__2172),
            .I(LED2_m0_rZ0));
    InMux I__433 (
            .O(N__2169),
            .I(N__2166));
    LocalMux I__432 (
            .O(N__2166),
            .I(N__2163));
    IoSpan4Mux I__431 (
            .O(N__2163),
            .I(N__2160));
    IoSpan4Mux I__430 (
            .O(N__2160),
            .I(N__2157));
    Odrv4 I__429 (
            .O(N__2157),
            .I(BUT2_c));
    CascadeMux I__428 (
            .O(N__2154),
            .I(N__2151));
    InMux I__427 (
            .O(N__2151),
            .I(N__2148));
    LocalMux I__426 (
            .O(N__2148),
            .I(N__2144));
    InMux I__425 (
            .O(N__2147),
            .I(N__2141));
    Span12Mux_s4_h I__424 (
            .O(N__2144),
            .I(N__2138));
    LocalMux I__423 (
            .O(N__2141),
            .I(BUT2_rZ0));
    Odrv12 I__422 (
            .O(N__2138),
            .I(BUT2_rZ0));
    InMux I__421 (
            .O(N__2133),
            .I(N__2128));
    InMux I__420 (
            .O(N__2132),
            .I(N__2125));
    InMux I__419 (
            .O(N__2131),
            .I(N__2122));
    LocalMux I__418 (
            .O(N__2128),
            .I(clk_divZ0Z_1));
    LocalMux I__417 (
            .O(N__2125),
            .I(clk_divZ0Z_1));
    LocalMux I__416 (
            .O(N__2122),
            .I(clk_divZ0Z_1));
    CascadeMux I__415 (
            .O(N__2115),
            .I(N__2109));
    CascadeMux I__414 (
            .O(N__2114),
            .I(N__2106));
    InMux I__413 (
            .O(N__2113),
            .I(N__2101));
    InMux I__412 (
            .O(N__2112),
            .I(N__2101));
    InMux I__411 (
            .O(N__2109),
            .I(N__2098));
    InMux I__410 (
            .O(N__2106),
            .I(N__2095));
    LocalMux I__409 (
            .O(N__2101),
            .I(clk_divZ0Z_0));
    LocalMux I__408 (
            .O(N__2098),
            .I(clk_divZ0Z_0));
    LocalMux I__407 (
            .O(N__2095),
            .I(clk_divZ0Z_0));
    CascadeMux I__406 (
            .O(N__2088),
            .I(N__2084));
    InMux I__405 (
            .O(N__2087),
            .I(N__2081));
    InMux I__404 (
            .O(N__2084),
            .I(N__2078));
    LocalMux I__403 (
            .O(N__2081),
            .I(clk_divZ0Z_2));
    LocalMux I__402 (
            .O(N__2078),
            .I(clk_divZ0Z_2));
    InMux I__401 (
            .O(N__2073),
            .I(clk_div_1_cry_1));
    CascadeMux I__400 (
            .O(N__2070),
            .I(N__2066));
    InMux I__399 (
            .O(N__2069),
            .I(N__2063));
    InMux I__398 (
            .O(N__2066),
            .I(N__2060));
    LocalMux I__397 (
            .O(N__2063),
            .I(clk_divZ0Z_3));
    LocalMux I__396 (
            .O(N__2060),
            .I(clk_divZ0Z_3));
    InMux I__395 (
            .O(N__2055),
            .I(clk_div_1_cry_2));
    CascadeMux I__394 (
            .O(N__2052),
            .I(N__2048));
    InMux I__393 (
            .O(N__2051),
            .I(N__2045));
    InMux I__392 (
            .O(N__2048),
            .I(N__2042));
    LocalMux I__391 (
            .O(N__2045),
            .I(clk_divZ0Z_4));
    LocalMux I__390 (
            .O(N__2042),
            .I(clk_divZ0Z_4));
    InMux I__389 (
            .O(N__2037),
            .I(clk_div_1_cry_3));
    InMux I__388 (
            .O(N__2034),
            .I(N__2031));
    LocalMux I__387 (
            .O(N__2031),
            .I(rst_cntZ0Z_13));
    InMux I__386 (
            .O(N__2028),
            .I(un1_rst_cnt_1_cry_12));
    InMux I__385 (
            .O(N__2025),
            .I(N__2021));
    InMux I__384 (
            .O(N__2024),
            .I(N__2018));
    LocalMux I__383 (
            .O(N__2021),
            .I(CONSTANT_ONE_NET));
    LocalMux I__382 (
            .O(N__2018),
            .I(CONSTANT_ONE_NET));
    InMux I__381 (
            .O(N__2013),
            .I(bfn_2_9_0_));
    InMux I__380 (
            .O(N__2010),
            .I(N__2005));
    InMux I__379 (
            .O(N__2009),
            .I(N__2000));
    InMux I__378 (
            .O(N__2008),
            .I(N__2000));
    LocalMux I__377 (
            .O(N__2005),
            .I(rst_cntZ0Z_14));
    LocalMux I__376 (
            .O(N__2000),
            .I(rst_cntZ0Z_14));
    CEMux I__375 (
            .O(N__1995),
            .I(N__1992));
    LocalMux I__374 (
            .O(N__1992),
            .I(N__1989));
    Span4Mux_h I__373 (
            .O(N__1989),
            .I(N__1986));
    Odrv4 I__372 (
            .O(N__1986),
            .I(N_16_0));
    SRMux I__371 (
            .O(N__1983),
            .I(N__1977));
    SRMux I__370 (
            .O(N__1982),
            .I(N__1974));
    SRMux I__369 (
            .O(N__1981),
            .I(N__1971));
    InMux I__368 (
            .O(N__1980),
            .I(N__1968));
    LocalMux I__367 (
            .O(N__1977),
            .I(BUT1_r_RNIKV9MZ0Z2));
    LocalMux I__366 (
            .O(N__1974),
            .I(BUT1_r_RNIKV9MZ0Z2));
    LocalMux I__365 (
            .O(N__1971),
            .I(BUT1_r_RNIKV9MZ0Z2));
    LocalMux I__364 (
            .O(N__1968),
            .I(BUT1_r_RNIKV9MZ0Z2));
    InMux I__363 (
            .O(N__1959),
            .I(N__1956));
    LocalMux I__362 (
            .O(N__1956),
            .I(N__1952));
    InMux I__361 (
            .O(N__1955),
            .I(N__1949));
    Odrv12 I__360 (
            .O(N__1952),
            .I(LED2_m1_rZ0));
    LocalMux I__359 (
            .O(N__1949),
            .I(LED2_m1_rZ0));
    IoInMux I__358 (
            .O(N__1944),
            .I(N__1941));
    LocalMux I__357 (
            .O(N__1941),
            .I(N__1938));
    Span4Mux_s3_h I__356 (
            .O(N__1938),
            .I(N__1935));
    Span4Mux_h I__355 (
            .O(N__1935),
            .I(N__1932));
    Odrv4 I__354 (
            .O(N__1932),
            .I(LED2_c));
    InMux I__353 (
            .O(N__1929),
            .I(N__1923));
    InMux I__352 (
            .O(N__1928),
            .I(N__1923));
    LocalMux I__351 (
            .O(N__1923),
            .I(N__1920));
    Span4Mux_h I__350 (
            .O(N__1920),
            .I(N__1917));
    Span4Mux_v I__349 (
            .O(N__1917),
            .I(N__1913));
    InMux I__348 (
            .O(N__1916),
            .I(N__1910));
    Odrv4 I__347 (
            .O(N__1913),
            .I(modeZ0));
    LocalMux I__346 (
            .O(N__1910),
            .I(modeZ0));
    InMux I__345 (
            .O(N__1905),
            .I(N__1902));
    LocalMux I__344 (
            .O(N__1902),
            .I(N__1898));
    InMux I__343 (
            .O(N__1901),
            .I(N__1895));
    Odrv4 I__342 (
            .O(N__1898),
            .I(LED1_m1_rZ0));
    LocalMux I__341 (
            .O(N__1895),
            .I(LED1_m1_rZ0));
    IoInMux I__340 (
            .O(N__1890),
            .I(N__1887));
    LocalMux I__339 (
            .O(N__1887),
            .I(N__1884));
    IoSpan4Mux I__338 (
            .O(N__1884),
            .I(N__1881));
    Span4Mux_s1_v I__337 (
            .O(N__1881),
            .I(N__1878));
    Odrv4 I__336 (
            .O(N__1878),
            .I(LED1_c));
    InMux I__335 (
            .O(N__1875),
            .I(N__1872));
    LocalMux I__334 (
            .O(N__1872),
            .I(rst_cntZ0Z_5));
    InMux I__333 (
            .O(N__1869),
            .I(un1_rst_cnt_1_cry_4));
    InMux I__332 (
            .O(N__1866),
            .I(N__1863));
    LocalMux I__331 (
            .O(N__1863),
            .I(rst_cntZ0Z_6));
    InMux I__330 (
            .O(N__1860),
            .I(un1_rst_cnt_1_cry_5));
    InMux I__329 (
            .O(N__1857),
            .I(N__1854));
    LocalMux I__328 (
            .O(N__1854),
            .I(rst_cntZ0Z_7));
    InMux I__327 (
            .O(N__1851),
            .I(un1_rst_cnt_1_cry_6));
    InMux I__326 (
            .O(N__1848),
            .I(N__1845));
    LocalMux I__325 (
            .O(N__1845),
            .I(rst_cntZ0Z_8));
    InMux I__324 (
            .O(N__1842),
            .I(bfn_2_8_0_));
    InMux I__323 (
            .O(N__1839),
            .I(N__1836));
    LocalMux I__322 (
            .O(N__1836),
            .I(rst_cntZ0Z_9));
    InMux I__321 (
            .O(N__1833),
            .I(un1_rst_cnt_1_cry_8));
    InMux I__320 (
            .O(N__1830),
            .I(N__1827));
    LocalMux I__319 (
            .O(N__1827),
            .I(rst_cntZ0Z_10));
    InMux I__318 (
            .O(N__1824),
            .I(un1_rst_cnt_1_cry_9));
    InMux I__317 (
            .O(N__1821),
            .I(N__1818));
    LocalMux I__316 (
            .O(N__1818),
            .I(rst_cntZ0Z_11));
    InMux I__315 (
            .O(N__1815),
            .I(un1_rst_cnt_1_cry_10));
    InMux I__314 (
            .O(N__1812),
            .I(N__1809));
    LocalMux I__313 (
            .O(N__1809),
            .I(rst_cntZ0Z_12));
    InMux I__312 (
            .O(N__1806),
            .I(un1_rst_cnt_1_cry_11));
    InMux I__311 (
            .O(N__1803),
            .I(N__1800));
    LocalMux I__310 (
            .O(N__1800),
            .I(cntr_1_9));
    CascadeMux I__309 (
            .O(N__1797),
            .I(N__1793));
    CascadeMux I__308 (
            .O(N__1796),
            .I(N__1790));
    InMux I__307 (
            .O(N__1793),
            .I(N__1784));
    InMux I__306 (
            .O(N__1790),
            .I(N__1784));
    InMux I__305 (
            .O(N__1789),
            .I(N__1781));
    LocalMux I__304 (
            .O(N__1784),
            .I(N__1778));
    LocalMux I__303 (
            .O(N__1781),
            .I(cntrZ0Z_9));
    Odrv4 I__302 (
            .O(N__1778),
            .I(cntrZ0Z_9));
    InMux I__301 (
            .O(N__1773),
            .I(N__1770));
    LocalMux I__300 (
            .O(N__1770),
            .I(cntr_1_11));
    InMux I__299 (
            .O(N__1767),
            .I(N__1762));
    InMux I__298 (
            .O(N__1766),
            .I(N__1759));
    InMux I__297 (
            .O(N__1765),
            .I(N__1756));
    LocalMux I__296 (
            .O(N__1762),
            .I(cntrZ0Z_11));
    LocalMux I__295 (
            .O(N__1759),
            .I(cntrZ0Z_11));
    LocalMux I__294 (
            .O(N__1756),
            .I(cntrZ0Z_11));
    CascadeMux I__293 (
            .O(N__1749),
            .I(N__1745));
    CascadeMux I__292 (
            .O(N__1748),
            .I(N__1738));
    InMux I__291 (
            .O(N__1745),
            .I(N__1730));
    InMux I__290 (
            .O(N__1744),
            .I(N__1725));
    InMux I__289 (
            .O(N__1743),
            .I(N__1725));
    InMux I__288 (
            .O(N__1742),
            .I(N__1722));
    CascadeMux I__287 (
            .O(N__1741),
            .I(N__1719));
    InMux I__286 (
            .O(N__1738),
            .I(N__1714));
    InMux I__285 (
            .O(N__1737),
            .I(N__1714));
    InMux I__284 (
            .O(N__1736),
            .I(N__1709));
    InMux I__283 (
            .O(N__1735),
            .I(N__1709));
    InMux I__282 (
            .O(N__1734),
            .I(N__1704));
    InMux I__281 (
            .O(N__1733),
            .I(N__1704));
    LocalMux I__280 (
            .O(N__1730),
            .I(N__1697));
    LocalMux I__279 (
            .O(N__1725),
            .I(N__1697));
    LocalMux I__278 (
            .O(N__1722),
            .I(N__1697));
    InMux I__277 (
            .O(N__1719),
            .I(N__1694));
    LocalMux I__276 (
            .O(N__1714),
            .I(cntrZ0Z_13));
    LocalMux I__275 (
            .O(N__1709),
            .I(cntrZ0Z_13));
    LocalMux I__274 (
            .O(N__1704),
            .I(cntrZ0Z_13));
    Odrv4 I__273 (
            .O(N__1697),
            .I(cntrZ0Z_13));
    LocalMux I__272 (
            .O(N__1694),
            .I(cntrZ0Z_13));
    InMux I__271 (
            .O(N__1683),
            .I(N__1680));
    LocalMux I__270 (
            .O(N__1680),
            .I(cntr_1_12));
    CascadeMux I__269 (
            .O(N__1677),
            .I(N__1672));
    CascadeMux I__268 (
            .O(N__1676),
            .I(N__1668));
    CascadeMux I__267 (
            .O(N__1675),
            .I(N__1665));
    InMux I__266 (
            .O(N__1672),
            .I(N__1655));
    InMux I__265 (
            .O(N__1671),
            .I(N__1655));
    InMux I__264 (
            .O(N__1668),
            .I(N__1655));
    InMux I__263 (
            .O(N__1665),
            .I(N__1652));
    CascadeMux I__262 (
            .O(N__1664),
            .I(N__1649));
    CascadeMux I__261 (
            .O(N__1663),
            .I(N__1646));
    CascadeMux I__260 (
            .O(N__1662),
            .I(N__1642));
    LocalMux I__259 (
            .O(N__1655),
            .I(N__1636));
    LocalMux I__258 (
            .O(N__1652),
            .I(N__1636));
    InMux I__257 (
            .O(N__1649),
            .I(N__1627));
    InMux I__256 (
            .O(N__1646),
            .I(N__1627));
    InMux I__255 (
            .O(N__1645),
            .I(N__1627));
    InMux I__254 (
            .O(N__1642),
            .I(N__1627));
    InMux I__253 (
            .O(N__1641),
            .I(N__1624));
    Span4Mux_s2_v I__252 (
            .O(N__1636),
            .I(N__1621));
    LocalMux I__251 (
            .O(N__1627),
            .I(cntrZ0Z_14));
    LocalMux I__250 (
            .O(N__1624),
            .I(cntrZ0Z_14));
    Odrv4 I__249 (
            .O(N__1621),
            .I(cntrZ0Z_14));
    CascadeMux I__248 (
            .O(N__1614),
            .I(N__1611));
    InMux I__247 (
            .O(N__1611),
            .I(N__1600));
    InMux I__246 (
            .O(N__1610),
            .I(N__1593));
    InMux I__245 (
            .O(N__1609),
            .I(N__1593));
    InMux I__244 (
            .O(N__1608),
            .I(N__1593));
    InMux I__243 (
            .O(N__1607),
            .I(N__1584));
    InMux I__242 (
            .O(N__1606),
            .I(N__1584));
    InMux I__241 (
            .O(N__1605),
            .I(N__1584));
    InMux I__240 (
            .O(N__1604),
            .I(N__1584));
    InMux I__239 (
            .O(N__1603),
            .I(N__1581));
    LocalMux I__238 (
            .O(N__1600),
            .I(cntr7lt13));
    LocalMux I__237 (
            .O(N__1593),
            .I(cntr7lt13));
    LocalMux I__236 (
            .O(N__1584),
            .I(cntr7lt13));
    LocalMux I__235 (
            .O(N__1581),
            .I(cntr7lt13));
    InMux I__234 (
            .O(N__1572),
            .I(N__1567));
    InMux I__233 (
            .O(N__1571),
            .I(N__1562));
    InMux I__232 (
            .O(N__1570),
            .I(N__1562));
    LocalMux I__231 (
            .O(N__1567),
            .I(cntrZ0Z_12));
    LocalMux I__230 (
            .O(N__1562),
            .I(cntrZ0Z_12));
    CascadeMux I__229 (
            .O(N__1557),
            .I(N__1553));
    InMux I__228 (
            .O(N__1556),
            .I(N__1550));
    InMux I__227 (
            .O(N__1553),
            .I(N__1547));
    LocalMux I__226 (
            .O(N__1550),
            .I(rst_cnt_i_14));
    LocalMux I__225 (
            .O(N__1547),
            .I(rst_cnt_i_14));
    InMux I__224 (
            .O(N__1542),
            .I(N__1539));
    LocalMux I__223 (
            .O(N__1539),
            .I(rst_cntZ0Z_0));
    InMux I__222 (
            .O(N__1536),
            .I(N__1533));
    LocalMux I__221 (
            .O(N__1533),
            .I(rst_cntZ0Z_1));
    InMux I__220 (
            .O(N__1530),
            .I(un1_rst_cnt_1_cry_0));
    InMux I__219 (
            .O(N__1527),
            .I(N__1524));
    LocalMux I__218 (
            .O(N__1524),
            .I(rst_cntZ0Z_2));
    InMux I__217 (
            .O(N__1521),
            .I(un1_rst_cnt_1_cry_1));
    InMux I__216 (
            .O(N__1518),
            .I(N__1515));
    LocalMux I__215 (
            .O(N__1515),
            .I(rst_cntZ0Z_3));
    InMux I__214 (
            .O(N__1512),
            .I(un1_rst_cnt_1_cry_2));
    InMux I__213 (
            .O(N__1509),
            .I(N__1506));
    LocalMux I__212 (
            .O(N__1506),
            .I(rst_cntZ0Z_4));
    InMux I__211 (
            .O(N__1503),
            .I(un1_rst_cnt_1_cry_3));
    CascadeMux I__210 (
            .O(N__1500),
            .I(cntr7lto7_0_4_cascade_));
    InMux I__209 (
            .O(N__1497),
            .I(N__1492));
    InMux I__208 (
            .O(N__1496),
            .I(N__1487));
    InMux I__207 (
            .O(N__1495),
            .I(N__1487));
    LocalMux I__206 (
            .O(N__1492),
            .I(cntrZ0Z_8));
    LocalMux I__205 (
            .O(N__1487),
            .I(cntrZ0Z_8));
    InMux I__204 (
            .O(N__1482),
            .I(N__1479));
    LocalMux I__203 (
            .O(N__1479),
            .I(LED1_m1_r_cnv_5));
    InMux I__202 (
            .O(N__1476),
            .I(N__1473));
    LocalMux I__201 (
            .O(N__1473),
            .I(N__1470));
    Odrv4 I__200 (
            .O(N__1470),
            .I(LED1_m1_r_cnv_6));
    InMux I__199 (
            .O(N__1467),
            .I(N__1464));
    LocalMux I__198 (
            .O(N__1464),
            .I(cntr7lto7_0_2));
    InMux I__197 (
            .O(N__1461),
            .I(N__1457));
    InMux I__196 (
            .O(N__1460),
            .I(N__1454));
    LocalMux I__195 (
            .O(N__1457),
            .I(N__1451));
    LocalMux I__194 (
            .O(N__1454),
            .I(cntrZ0Z_2));
    Odrv4 I__193 (
            .O(N__1451),
            .I(cntrZ0Z_2));
    CascadeMux I__192 (
            .O(N__1446),
            .I(N__1442));
    InMux I__191 (
            .O(N__1445),
            .I(N__1439));
    InMux I__190 (
            .O(N__1442),
            .I(N__1436));
    LocalMux I__189 (
            .O(N__1439),
            .I(cntrZ0Z_3));
    LocalMux I__188 (
            .O(N__1436),
            .I(cntrZ0Z_3));
    InMux I__187 (
            .O(N__1431),
            .I(N__1427));
    InMux I__186 (
            .O(N__1430),
            .I(N__1424));
    LocalMux I__185 (
            .O(N__1427),
            .I(cntr7lt5_3));
    LocalMux I__184 (
            .O(N__1424),
            .I(cntr7lt5_3));
    InMux I__183 (
            .O(N__1419),
            .I(N__1414));
    InMux I__182 (
            .O(N__1418),
            .I(N__1409));
    InMux I__181 (
            .O(N__1417),
            .I(N__1409));
    LocalMux I__180 (
            .O(N__1414),
            .I(cntrZ0Z_6));
    LocalMux I__179 (
            .O(N__1409),
            .I(cntrZ0Z_6));
    InMux I__178 (
            .O(N__1404),
            .I(N__1398));
    InMux I__177 (
            .O(N__1403),
            .I(N__1395));
    InMux I__176 (
            .O(N__1402),
            .I(N__1390));
    InMux I__175 (
            .O(N__1401),
            .I(N__1390));
    LocalMux I__174 (
            .O(N__1398),
            .I(cntrZ0Z_5));
    LocalMux I__173 (
            .O(N__1395),
            .I(cntrZ0Z_5));
    LocalMux I__172 (
            .O(N__1390),
            .I(cntrZ0Z_5));
    CascadeMux I__171 (
            .O(N__1383),
            .I(N__1379));
    InMux I__170 (
            .O(N__1382),
            .I(N__1372));
    InMux I__169 (
            .O(N__1379),
            .I(N__1372));
    InMux I__168 (
            .O(N__1378),
            .I(N__1369));
    InMux I__167 (
            .O(N__1377),
            .I(N__1366));
    LocalMux I__166 (
            .O(N__1372),
            .I(N__1363));
    LocalMux I__165 (
            .O(N__1369),
            .I(cntrZ0Z_7));
    LocalMux I__164 (
            .O(N__1366),
            .I(cntrZ0Z_7));
    Odrv4 I__163 (
            .O(N__1363),
            .I(cntrZ0Z_7));
    InMux I__162 (
            .O(N__1356),
            .I(N__1351));
    InMux I__161 (
            .O(N__1355),
            .I(N__1346));
    InMux I__160 (
            .O(N__1354),
            .I(N__1346));
    LocalMux I__159 (
            .O(N__1351),
            .I(cntrZ0Z_4));
    LocalMux I__158 (
            .O(N__1346),
            .I(cntrZ0Z_4));
    InMux I__157 (
            .O(N__1341),
            .I(N__1338));
    LocalMux I__156 (
            .O(N__1338),
            .I(cntr7lto7_c));
    InMux I__155 (
            .O(N__1335),
            .I(N__1332));
    LocalMux I__154 (
            .O(N__1332),
            .I(cntr_1_10));
    InMux I__153 (
            .O(N__1329),
            .I(N__1324));
    InMux I__152 (
            .O(N__1328),
            .I(N__1319));
    InMux I__151 (
            .O(N__1327),
            .I(N__1319));
    LocalMux I__150 (
            .O(N__1324),
            .I(cntrZ0Z_10));
    LocalMux I__149 (
            .O(N__1319),
            .I(cntrZ0Z_10));
    InMux I__148 (
            .O(N__1314),
            .I(N__1306));
    InMux I__147 (
            .O(N__1313),
            .I(N__1306));
    InMux I__146 (
            .O(N__1312),
            .I(N__1303));
    InMux I__145 (
            .O(N__1311),
            .I(N__1300));
    LocalMux I__144 (
            .O(N__1306),
            .I(cntrZ0Z_0));
    LocalMux I__143 (
            .O(N__1303),
            .I(cntrZ0Z_0));
    LocalMux I__142 (
            .O(N__1300),
            .I(cntrZ0Z_0));
    CascadeMux I__141 (
            .O(N__1293),
            .I(N__1289));
    InMux I__140 (
            .O(N__1292),
            .I(N__1285));
    InMux I__139 (
            .O(N__1289),
            .I(N__1282));
    InMux I__138 (
            .O(N__1288),
            .I(N__1279));
    LocalMux I__137 (
            .O(N__1285),
            .I(cntrZ0Z_1));
    LocalMux I__136 (
            .O(N__1282),
            .I(cntrZ0Z_1));
    LocalMux I__135 (
            .O(N__1279),
            .I(cntrZ0Z_1));
    CascadeMux I__134 (
            .O(N__1272),
            .I(BUT1_r_RNIKV9MZ0Z2_cascade_));
    SRMux I__133 (
            .O(N__1269),
            .I(N__1266));
    LocalMux I__132 (
            .O(N__1266),
            .I(N__1263));
    Odrv12 I__131 (
            .O(N__1263),
            .I(cntr_RNITQ4V2Z0Z_14));
    CascadeMux I__130 (
            .O(N__1260),
            .I(LED1_m1_r_cnv_7_cascade_));
    InMux I__129 (
            .O(N__1257),
            .I(N__1251));
    InMux I__128 (
            .O(N__1256),
            .I(N__1251));
    LocalMux I__127 (
            .O(N__1251),
            .I(cntr_RNIV9NN2Z0Z_4));
    InMux I__126 (
            .O(N__1248),
            .I(bfn_1_5_0_));
    InMux I__125 (
            .O(N__1245),
            .I(cntr_1_cry_9));
    InMux I__124 (
            .O(N__1242),
            .I(cntr_1_cry_10));
    InMux I__123 (
            .O(N__1239),
            .I(cntr_1_cry_11));
    InMux I__122 (
            .O(N__1236),
            .I(cntr_1_cry_12));
    InMux I__121 (
            .O(N__1233),
            .I(cntr_1_cry_13));
    IoInMux I__120 (
            .O(N__1230),
            .I(N__1227));
    LocalMux I__119 (
            .O(N__1227),
            .I(clk_div_RNIM1KP1Z0Z_11));
    InMux I__118 (
            .O(N__1224),
            .I(cntr_1_cry_1));
    InMux I__117 (
            .O(N__1221),
            .I(cntr_1_cry_2));
    InMux I__116 (
            .O(N__1218),
            .I(cntr_1_cry_3));
    InMux I__115 (
            .O(N__1215),
            .I(N__1212));
    LocalMux I__114 (
            .O(N__1212),
            .I(cntr_1_5));
    InMux I__113 (
            .O(N__1209),
            .I(cntr_1_cry_4));
    InMux I__112 (
            .O(N__1206),
            .I(N__1203));
    LocalMux I__111 (
            .O(N__1203),
            .I(cntr_1_6));
    InMux I__110 (
            .O(N__1200),
            .I(cntr_1_cry_5));
    InMux I__109 (
            .O(N__1197),
            .I(cntr_1_cry_6));
    InMux I__108 (
            .O(N__1194),
            .I(N__1191));
    LocalMux I__107 (
            .O(N__1191),
            .I(cntr_1_8));
    InMux I__106 (
            .O(N__1188),
            .I(cntr_1_cry_7));
    defparam IN_MUX_bfv_1_4_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_4_0_ (
            .carryinitin(),
            .carryinitout(bfn_1_4_0_));
    defparam IN_MUX_bfv_1_5_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_1_5_0_ (
            .carryinitin(cntr_1_cry_8),
            .carryinitout(bfn_1_5_0_));
    defparam IN_MUX_bfv_4_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_4_7_0_));
    defparam IN_MUX_bfv_4_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_4_8_0_ (
            .carryinitin(clk_div_2_cry_8),
            .carryinitout(bfn_4_8_0_));
    defparam IN_MUX_bfv_5_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_5_7_0_));
    defparam IN_MUX_bfv_5_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_5_8_0_ (
            .carryinitin(clk_div_1_cry_8),
            .carryinitout(bfn_5_8_0_));
    defparam IN_MUX_bfv_2_7_0_.C_INIT=2'b00;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_7_0_ (
            .carryinitin(),
            .carryinitout(bfn_2_7_0_));
    defparam IN_MUX_bfv_2_8_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_8_0_ (
            .carryinitin(un1_rst_cnt_1_cry_7),
            .carryinitout(bfn_2_8_0_));
    defparam IN_MUX_bfv_2_9_0_.C_INIT=2'b10;
    ICE_CARRY_IN_MUX IN_MUX_bfv_2_9_0_ (
            .carryinitin(un1_rst_cnt_1_cry_13_THRU_CRY_1_THRU_CO),
            .carryinitout(bfn_2_9_0_));
    VCC VCC (
            .Y(VCCG0));
    GND GND (
            .Y(GNDG0));
    ICE_GB clk_div_RNIM1KP1_0_11 (
            .USERSIGNALTOGLOBALBUFFER(N__1230),
            .GLOBALBUFFEROUTPUT(N_16_g));
    GND GND_Inst (
            .Y(_gnd_net_));
    defparam cntr_5_LC_1_3_3.C_ON=1'b0;
    defparam cntr_5_LC_1_3_3.SEQ_MODE=4'b1000;
    defparam cntr_5_LC_1_3_3.LUT_INIT=16'b0000110001001100;
    LogicCell40 cntr_5_LC_1_3_3 (
            .in0(N__1743),
            .in1(N__1215),
            .in2(N__1676),
            .in3(N__1609),
            .lcout(cntrZ0Z_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2377),
            .ce(N__2269),
            .sr(_gnd_net_));
    defparam cntr_6_LC_1_3_6.C_ON=1'b0;
    defparam cntr_6_LC_1_3_6.SEQ_MODE=4'b1000;
    defparam cntr_6_LC_1_3_6.LUT_INIT=16'b0011011100000000;
    LogicCell40 cntr_6_LC_1_3_6 (
            .in0(N__1608),
            .in1(N__1671),
            .in2(N__1749),
            .in3(N__1206),
            .lcout(cntrZ0Z_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2377),
            .ce(N__2269),
            .sr(_gnd_net_));
    defparam cntr_8_LC_1_3_7.C_ON=1'b0;
    defparam cntr_8_LC_1_3_7.SEQ_MODE=4'b1000;
    defparam cntr_8_LC_1_3_7.LUT_INIT=16'b0000110001001100;
    LogicCell40 cntr_8_LC_1_3_7 (
            .in0(N__1744),
            .in1(N__1194),
            .in2(N__1677),
            .in3(N__1610),
            .lcout(cntrZ0Z_8),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2377),
            .ce(N__2269),
            .sr(_gnd_net_));
    defparam cntr_1_cry_1_c_LC_1_4_0.C_ON=1'b1;
    defparam cntr_1_cry_1_c_LC_1_4_0.SEQ_MODE=4'b0000;
    defparam cntr_1_cry_1_c_LC_1_4_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 cntr_1_cry_1_c_LC_1_4_0 (
            .in0(_gnd_net_),
            .in1(N__1312),
            .in2(N__1293),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_1_4_0_),
            .carryout(cntr_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_2_LC_1_4_1.C_ON=1'b1;
    defparam cntr_2_LC_1_4_1.SEQ_MODE=4'b1000;
    defparam cntr_2_LC_1_4_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntr_2_LC_1_4_1 (
            .in0(_gnd_net_),
            .in1(N__1460),
            .in2(_gnd_net_),
            .in3(N__1224),
            .lcout(cntrZ0Z_2),
            .ltout(),
            .carryin(cntr_1_cry_1),
            .carryout(cntr_1_cry_2),
            .clk(N__2375),
            .ce(N__2267),
            .sr(_gnd_net_));
    defparam cntr_3_LC_1_4_2.C_ON=1'b1;
    defparam cntr_3_LC_1_4_2.SEQ_MODE=4'b1000;
    defparam cntr_3_LC_1_4_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntr_3_LC_1_4_2 (
            .in0(_gnd_net_),
            .in1(N__1445),
            .in2(_gnd_net_),
            .in3(N__1221),
            .lcout(cntrZ0Z_3),
            .ltout(),
            .carryin(cntr_1_cry_2),
            .carryout(cntr_1_cry_3),
            .clk(N__2375),
            .ce(N__2267),
            .sr(_gnd_net_));
    defparam cntr_4_LC_1_4_3.C_ON=1'b1;
    defparam cntr_4_LC_1_4_3.SEQ_MODE=4'b1000;
    defparam cntr_4_LC_1_4_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntr_4_LC_1_4_3 (
            .in0(_gnd_net_),
            .in1(N__1356),
            .in2(_gnd_net_),
            .in3(N__1218),
            .lcout(cntrZ0Z_4),
            .ltout(),
            .carryin(cntr_1_cry_3),
            .carryout(cntr_1_cry_4),
            .clk(N__2375),
            .ce(N__2267),
            .sr(_gnd_net_));
    defparam cntr_RNO_0_5_LC_1_4_4.C_ON=1'b1;
    defparam cntr_RNO_0_5_LC_1_4_4.SEQ_MODE=4'b0000;
    defparam cntr_RNO_0_5_LC_1_4_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntr_RNO_0_5_LC_1_4_4 (
            .in0(_gnd_net_),
            .in1(N__1403),
            .in2(_gnd_net_),
            .in3(N__1209),
            .lcout(cntr_1_5),
            .ltout(),
            .carryin(cntr_1_cry_4),
            .carryout(cntr_1_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNO_0_6_LC_1_4_5.C_ON=1'b1;
    defparam cntr_RNO_0_6_LC_1_4_5.SEQ_MODE=4'b0000;
    defparam cntr_RNO_0_6_LC_1_4_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntr_RNO_0_6_LC_1_4_5 (
            .in0(_gnd_net_),
            .in1(N__1419),
            .in2(_gnd_net_),
            .in3(N__1200),
            .lcout(cntr_1_6),
            .ltout(),
            .carryin(cntr_1_cry_5),
            .carryout(cntr_1_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_7_LC_1_4_6.C_ON=1'b1;
    defparam cntr_7_LC_1_4_6.SEQ_MODE=4'b1000;
    defparam cntr_7_LC_1_4_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntr_7_LC_1_4_6 (
            .in0(_gnd_net_),
            .in1(N__1377),
            .in2(_gnd_net_),
            .in3(N__1197),
            .lcout(cntrZ0Z_7),
            .ltout(),
            .carryin(cntr_1_cry_6),
            .carryout(cntr_1_cry_7),
            .clk(N__2375),
            .ce(N__2267),
            .sr(_gnd_net_));
    defparam cntr_RNO_0_8_LC_1_4_7.C_ON=1'b1;
    defparam cntr_RNO_0_8_LC_1_4_7.SEQ_MODE=4'b0000;
    defparam cntr_RNO_0_8_LC_1_4_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntr_RNO_0_8_LC_1_4_7 (
            .in0(_gnd_net_),
            .in1(N__1497),
            .in2(_gnd_net_),
            .in3(N__1188),
            .lcout(cntr_1_8),
            .ltout(),
            .carryin(cntr_1_cry_7),
            .carryout(cntr_1_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNO_0_9_LC_1_5_0.C_ON=1'b1;
    defparam cntr_RNO_0_9_LC_1_5_0.SEQ_MODE=4'b0000;
    defparam cntr_RNO_0_9_LC_1_5_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntr_RNO_0_9_LC_1_5_0 (
            .in0(_gnd_net_),
            .in1(N__1789),
            .in2(_gnd_net_),
            .in3(N__1248),
            .lcout(cntr_1_9),
            .ltout(),
            .carryin(bfn_1_5_0_),
            .carryout(cntr_1_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNO_0_10_LC_1_5_1.C_ON=1'b1;
    defparam cntr_RNO_0_10_LC_1_5_1.SEQ_MODE=4'b0000;
    defparam cntr_RNO_0_10_LC_1_5_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntr_RNO_0_10_LC_1_5_1 (
            .in0(_gnd_net_),
            .in1(N__1329),
            .in2(_gnd_net_),
            .in3(N__1245),
            .lcout(cntr_1_10),
            .ltout(),
            .carryin(cntr_1_cry_9),
            .carryout(cntr_1_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNO_0_11_LC_1_5_2.C_ON=1'b1;
    defparam cntr_RNO_0_11_LC_1_5_2.SEQ_MODE=4'b0000;
    defparam cntr_RNO_0_11_LC_1_5_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntr_RNO_0_11_LC_1_5_2 (
            .in0(_gnd_net_),
            .in1(N__1767),
            .in2(_gnd_net_),
            .in3(N__1242),
            .lcout(cntr_1_11),
            .ltout(),
            .carryin(cntr_1_cry_10),
            .carryout(cntr_1_cry_11),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNO_0_12_LC_1_5_3.C_ON=1'b1;
    defparam cntr_RNO_0_12_LC_1_5_3.SEQ_MODE=4'b0000;
    defparam cntr_RNO_0_12_LC_1_5_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntr_RNO_0_12_LC_1_5_3 (
            .in0(_gnd_net_),
            .in1(N__1572),
            .in2(_gnd_net_),
            .in3(N__1239),
            .lcout(cntr_1_12),
            .ltout(),
            .carryin(cntr_1_cry_11),
            .carryout(cntr_1_cry_12),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_13_LC_1_5_4.C_ON=1'b1;
    defparam cntr_13_LC_1_5_4.SEQ_MODE=4'b1000;
    defparam cntr_13_LC_1_5_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 cntr_13_LC_1_5_4 (
            .in0(_gnd_net_),
            .in1(N__1733),
            .in2(_gnd_net_),
            .in3(N__1236),
            .lcout(cntrZ0Z_13),
            .ltout(),
            .carryin(cntr_1_cry_12),
            .carryout(cntr_1_cry_13),
            .clk(N__2373),
            .ce(N__2266),
            .sr(_gnd_net_));
    defparam cntr_14_LC_1_5_5.C_ON=1'b0;
    defparam cntr_14_LC_1_5_5.SEQ_MODE=4'b1000;
    defparam cntr_14_LC_1_5_5.LUT_INIT=16'b0011001100000100;
    LogicCell40 cntr_14_LC_1_5_5 (
            .in0(N__1734),
            .in1(N__1641),
            .in2(N__1614),
            .in3(N__1233),
            .lcout(cntrZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2373),
            .ce(N__2266),
            .sr(_gnd_net_));
    defparam mode_LC_1_7_3.C_ON=1'b0;
    defparam mode_LC_1_7_3.SEQ_MODE=4'b1000;
    defparam mode_LC_1_7_3.LUT_INIT=16'b0011001111001100;
    LogicCell40 mode_LC_1_7_3 (
            .in0(_gnd_net_),
            .in1(N__1916),
            .in2(_gnd_net_),
            .in3(N__1980),
            .lcout(modeZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2369),
            .ce(),
            .sr(_gnd_net_));
    defparam CONSTANT_ONE_LUT4_LC_1_8_0.C_ON=1'b0;
    defparam CONSTANT_ONE_LUT4_LC_1_8_0.SEQ_MODE=4'b0000;
    defparam CONSTANT_ONE_LUT4_LC_1_8_0.LUT_INIT=16'b1111111111111111;
    LogicCell40 CONSTANT_ONE_LUT4_LC_1_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(CONSTANT_ONE_NET),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNIM1KP1_11_LC_1_8_2.C_ON=1'b0;
    defparam clk_div_RNIM1KP1_11_LC_1_8_2.SEQ_MODE=4'b0000;
    defparam clk_div_RNIM1KP1_11_LC_1_8_2.LUT_INIT=16'b0000000011110000;
    LogicCell40 clk_div_RNIM1KP1_11_LC_1_8_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2214),
            .in3(N__2196),
            .lcout(clk_div_RNIM1KP1Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rst_cnt_esr_RNI37G6_14_LC_1_8_3.C_ON=1'b0;
    defparam rst_cnt_esr_RNI37G6_14_LC_1_8_3.SEQ_MODE=4'b0000;
    defparam rst_cnt_esr_RNI37G6_14_LC_1_8_3.LUT_INIT=16'b0000000011111111;
    LogicCell40 rst_cnt_esr_RNI37G6_14_LC_1_8_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2008),
            .lcout(rst_cnt_i_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam BUT1_r_RNIKV9M2_LC_1_8_5.C_ON=1'b0;
    defparam BUT1_r_RNIKV9M2_LC_1_8_5.SEQ_MODE=4'b0000;
    defparam BUT1_r_RNIKV9M2_LC_1_8_5.LUT_INIT=16'b0000010000000000;
    LogicCell40 BUT1_r_RNIKV9M2_LC_1_8_5 (
            .in0(N__2403),
            .in1(N__2009),
            .in2(N__2154),
            .in3(N__2314),
            .lcout(BUT1_r_RNIKV9MZ0Z2),
            .ltout(BUT1_r_RNIKV9MZ0Z2_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rst_cnt_esr_RNO_0_14_LC_1_8_6.C_ON=1'b0;
    defparam rst_cnt_esr_RNO_0_14_LC_1_8_6.SEQ_MODE=4'b0000;
    defparam rst_cnt_esr_RNO_0_14_LC_1_8_6.LUT_INIT=16'b1111101011111010;
    LogicCell40 rst_cnt_esr_RNO_0_14_LC_1_8_6 (
            .in0(N__2315),
            .in1(_gnd_net_),
            .in2(N__1272),
            .in3(_gnd_net_),
            .lcout(N_16_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LED1_m1_r_LC_2_2_3.C_ON=1'b0;
    defparam LED1_m1_r_LC_2_2_3.SEQ_MODE=4'b1001;
    defparam LED1_m1_r_LC_2_2_3.LUT_INIT=16'b0000000011001100;
    LogicCell40 LED1_m1_r_LC_2_2_3 (
            .in0(_gnd_net_),
            .in1(N__1901),
            .in2(_gnd_net_),
            .in3(N__1256),
            .lcout(LED1_m1_rZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2380),
            .ce(),
            .sr(N__1269));
    defparam LED2_m1_r_LC_2_2_5.C_ON=1'b0;
    defparam LED2_m1_r_LC_2_2_5.SEQ_MODE=4'b1000;
    defparam LED2_m1_r_LC_2_2_5.LUT_INIT=16'b1111111110101010;
    LogicCell40 LED2_m1_r_LC_2_2_5 (
            .in0(N__1955),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1257),
            .lcout(LED2_m1_rZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2380),
            .ce(),
            .sr(N__1269));
    defparam cntr_RNITQ4V2_14_LC_2_3_1.C_ON=1'b0;
    defparam cntr_RNITQ4V2_14_LC_2_3_1.SEQ_MODE=4'b0000;
    defparam cntr_RNITQ4V2_14_LC_2_3_1.LUT_INIT=16'b1110000000000000;
    LogicCell40 cntr_RNITQ4V2_14_LC_2_3_1 (
            .in0(N__1742),
            .in1(N__1603),
            .in2(N__1675),
            .in3(N__2316),
            .lcout(cntr_RNITQ4V2Z0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNIGH28_5_LC_2_3_4.C_ON=1'b0;
    defparam cntr_RNIGH28_5_LC_2_3_4.SEQ_MODE=4'b0000;
    defparam cntr_RNIGH28_5_LC_2_3_4.LUT_INIT=16'b1000100000000000;
    LogicCell40 cntr_RNIGH28_5_LC_2_3_4 (
            .in0(N__1482),
            .in1(N__1378),
            .in2(_gnd_net_),
            .in3(N__1404),
            .lcout(),
            .ltout(LED1_m1_r_cnv_7_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNIV9NN2_4_LC_2_3_5.C_ON=1'b0;
    defparam cntr_RNIV9NN2_4_LC_2_3_5.SEQ_MODE=4'b0000;
    defparam cntr_RNIV9NN2_4_LC_2_3_5.LUT_INIT=16'b1000000000000000;
    LogicCell40 cntr_RNIV9NN2_4_LC_2_3_5 (
            .in0(N__1476),
            .in1(N__1431),
            .in2(N__1260),
            .in3(N__2317),
            .lcout(cntr_RNIV9NN2Z0Z_4),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNIKC8M_8_LC_2_4_0.C_ON=1'b0;
    defparam cntr_RNIKC8M_8_LC_2_4_0.SEQ_MODE=4'b0000;
    defparam cntr_RNIKC8M_8_LC_2_4_0.LUT_INIT=16'b1000000000000000;
    LogicCell40 cntr_RNIKC8M_8_LC_2_4_0 (
            .in0(N__1496),
            .in1(N__1341),
            .in2(N__1797),
            .in3(N__1467),
            .lcout(),
            .ltout(cntr7lto7_0_4_cascade_),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNI0LHN_5_LC_2_4_1.C_ON=1'b0;
    defparam cntr_RNI0LHN_5_LC_2_4_1.SEQ_MODE=4'b0000;
    defparam cntr_RNI0LHN_5_LC_2_4_1.LUT_INIT=16'b1111000011100000;
    LogicCell40 cntr_RNI0LHN_5_LC_2_4_1 (
            .in0(N__1382),
            .in1(N__1430),
            .in2(N__1500),
            .in3(N__1402),
            .lcout(cntr7lt13),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNI6JK7_6_LC_2_4_2.C_ON=1'b0;
    defparam cntr_RNI6JK7_6_LC_2_4_2.SEQ_MODE=4'b0000;
    defparam cntr_RNI6JK7_6_LC_2_4_2.LUT_INIT=16'b0000000000100000;
    LogicCell40 cntr_RNI6JK7_6_LC_2_4_2 (
            .in0(N__1495),
            .in1(N__1418),
            .in2(N__1796),
            .in3(N__1571),
            .lcout(LED1_m1_r_cnv_5),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNINC5L_4_LC_2_4_3.C_ON=1'b0;
    defparam cntr_RNINC5L_4_LC_2_4_3.SEQ_MODE=4'b0000;
    defparam cntr_RNINC5L_4_LC_2_4_3.LUT_INIT=16'b0010000000000000;
    LogicCell40 cntr_RNINC5L_4_LC_2_4_3 (
            .in0(N__1766),
            .in1(N__1355),
            .in2(N__1741),
            .in3(N__1328),
            .lcout(LED1_m1_r_cnv_6),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNIJEUK_10_LC_2_4_5.C_ON=1'b0;
    defparam cntr_RNIJEUK_10_LC_2_4_5.SEQ_MODE=4'b0000;
    defparam cntr_RNIJEUK_10_LC_2_4_5.LUT_INIT=16'b1000100000000000;
    LogicCell40 cntr_RNIJEUK_10_LC_2_4_5 (
            .in0(N__1570),
            .in1(N__1765),
            .in2(_gnd_net_),
            .in3(N__1327),
            .lcout(cntr7lto7_0_2),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNI2AR_1_LC_2_4_6.C_ON=1'b0;
    defparam cntr_RNI2AR_1_LC_2_4_6.SEQ_MODE=4'b0000;
    defparam cntr_RNI2AR_1_LC_2_4_6.LUT_INIT=16'b1000000000000000;
    LogicCell40 cntr_RNI2AR_1_LC_2_4_6 (
            .in0(N__1461),
            .in1(N__1288),
            .in2(N__1446),
            .in3(N__1311),
            .lcout(cntr7lt5_3),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_RNIIQR_4_LC_2_4_7.C_ON=1'b0;
    defparam cntr_RNIIQR_4_LC_2_4_7.SEQ_MODE=4'b0000;
    defparam cntr_RNIIQR_4_LC_2_4_7.LUT_INIT=16'b1111101011111000;
    LogicCell40 cntr_RNIIQR_4_LC_2_4_7 (
            .in0(N__1417),
            .in1(N__1401),
            .in2(N__1383),
            .in3(N__1354),
            .lcout(cntr7lto7_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam cntr_0_LC_2_5_0.C_ON=1'b0;
    defparam cntr_0_LC_2_5_0.SEQ_MODE=4'b1000;
    defparam cntr_0_LC_2_5_0.LUT_INIT=16'b0000000011111111;
    LogicCell40 cntr_0_LC_2_5_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__1313),
            .lcout(cntrZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2376),
            .ce(N__2268),
            .sr(_gnd_net_));
    defparam cntr_10_LC_2_5_1.C_ON=1'b0;
    defparam cntr_10_LC_2_5_1.SEQ_MODE=4'b1000;
    defparam cntr_10_LC_2_5_1.LUT_INIT=16'b0000101000101010;
    LogicCell40 cntr_10_LC_2_5_1 (
            .in0(N__1335),
            .in1(N__1737),
            .in2(N__1662),
            .in3(N__1605),
            .lcout(cntrZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2376),
            .ce(N__2268),
            .sr(_gnd_net_));
    defparam cntr_1_LC_2_5_2.C_ON=1'b0;
    defparam cntr_1_LC_2_5_2.SEQ_MODE=4'b1000;
    defparam cntr_1_LC_2_5_2.LUT_INIT=16'b1100001100111100;
    LogicCell40 cntr_1_LC_2_5_2 (
            .in0(_gnd_net_),
            .in1(N__1292),
            .in2(_gnd_net_),
            .in3(N__1314),
            .lcout(cntrZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2376),
            .ce(N__2268),
            .sr(_gnd_net_));
    defparam cntr_9_LC_2_5_3.C_ON=1'b0;
    defparam cntr_9_LC_2_5_3.SEQ_MODE=4'b1000;
    defparam cntr_9_LC_2_5_3.LUT_INIT=16'b0000110001001100;
    LogicCell40 cntr_9_LC_2_5_3 (
            .in0(N__1736),
            .in1(N__1803),
            .in2(N__1664),
            .in3(N__1607),
            .lcout(cntrZ0Z_9),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2376),
            .ce(N__2268),
            .sr(_gnd_net_));
    defparam cntr_11_LC_2_5_6.C_ON=1'b0;
    defparam cntr_11_LC_2_5_6.SEQ_MODE=4'b1000;
    defparam cntr_11_LC_2_5_6.LUT_INIT=16'b0011011100000000;
    LogicCell40 cntr_11_LC_2_5_6 (
            .in0(N__1604),
            .in1(N__1645),
            .in2(N__1748),
            .in3(N__1773),
            .lcout(cntrZ0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2376),
            .ce(N__2268),
            .sr(_gnd_net_));
    defparam cntr_12_LC_2_5_7.C_ON=1'b0;
    defparam cntr_12_LC_2_5_7.SEQ_MODE=4'b1000;
    defparam cntr_12_LC_2_5_7.LUT_INIT=16'b0000110001001100;
    LogicCell40 cntr_12_LC_2_5_7 (
            .in0(N__1735),
            .in1(N__1683),
            .in2(N__1663),
            .in3(N__1606),
            .lcout(cntrZ0Z_12),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2376),
            .ce(N__2268),
            .sr(_gnd_net_));
    defparam rst_cnt_0_LC_2_7_0.C_ON=1'b1;
    defparam rst_cnt_0_LC_2_7_0.SEQ_MODE=4'b1000;
    defparam rst_cnt_0_LC_2_7_0.LUT_INIT=16'b0110011011001100;
    LogicCell40 rst_cnt_0_LC_2_7_0 (
            .in0(N__2328),
            .in1(N__1542),
            .in2(N__1557),
            .in3(N__1556),
            .lcout(rst_cntZ0Z_0),
            .ltout(),
            .carryin(bfn_2_7_0_),
            .carryout(un1_rst_cnt_1_cry_0),
            .clk(N__2370),
            .ce(),
            .sr(N__1982));
    defparam rst_cnt_1_LC_2_7_1.C_ON=1'b1;
    defparam rst_cnt_1_LC_2_7_1.SEQ_MODE=4'b1000;
    defparam rst_cnt_1_LC_2_7_1.LUT_INIT=16'b0110011011001100;
    LogicCell40 rst_cnt_1_LC_2_7_1 (
            .in0(N__2321),
            .in1(N__1536),
            .in2(_gnd_net_),
            .in3(N__1530),
            .lcout(rst_cntZ0Z_1),
            .ltout(),
            .carryin(un1_rst_cnt_1_cry_0),
            .carryout(un1_rst_cnt_1_cry_1),
            .clk(N__2370),
            .ce(),
            .sr(N__1982));
    defparam rst_cnt_2_LC_2_7_2.C_ON=1'b1;
    defparam rst_cnt_2_LC_2_7_2.SEQ_MODE=4'b1000;
    defparam rst_cnt_2_LC_2_7_2.LUT_INIT=16'b0110011011001100;
    LogicCell40 rst_cnt_2_LC_2_7_2 (
            .in0(N__2329),
            .in1(N__1527),
            .in2(_gnd_net_),
            .in3(N__1521),
            .lcout(rst_cntZ0Z_2),
            .ltout(),
            .carryin(un1_rst_cnt_1_cry_1),
            .carryout(un1_rst_cnt_1_cry_2),
            .clk(N__2370),
            .ce(),
            .sr(N__1982));
    defparam rst_cnt_3_LC_2_7_3.C_ON=1'b1;
    defparam rst_cnt_3_LC_2_7_3.SEQ_MODE=4'b1000;
    defparam rst_cnt_3_LC_2_7_3.LUT_INIT=16'b0110011011001100;
    LogicCell40 rst_cnt_3_LC_2_7_3 (
            .in0(N__2322),
            .in1(N__1518),
            .in2(_gnd_net_),
            .in3(N__1512),
            .lcout(rst_cntZ0Z_3),
            .ltout(),
            .carryin(un1_rst_cnt_1_cry_2),
            .carryout(un1_rst_cnt_1_cry_3),
            .clk(N__2370),
            .ce(),
            .sr(N__1982));
    defparam rst_cnt_4_LC_2_7_4.C_ON=1'b1;
    defparam rst_cnt_4_LC_2_7_4.SEQ_MODE=4'b1000;
    defparam rst_cnt_4_LC_2_7_4.LUT_INIT=16'b0110011011001100;
    LogicCell40 rst_cnt_4_LC_2_7_4 (
            .in0(N__2330),
            .in1(N__1509),
            .in2(_gnd_net_),
            .in3(N__1503),
            .lcout(rst_cntZ0Z_4),
            .ltout(),
            .carryin(un1_rst_cnt_1_cry_3),
            .carryout(un1_rst_cnt_1_cry_4),
            .clk(N__2370),
            .ce(),
            .sr(N__1982));
    defparam rst_cnt_5_LC_2_7_5.C_ON=1'b1;
    defparam rst_cnt_5_LC_2_7_5.SEQ_MODE=4'b1000;
    defparam rst_cnt_5_LC_2_7_5.LUT_INIT=16'b0110011011001100;
    LogicCell40 rst_cnt_5_LC_2_7_5 (
            .in0(N__2323),
            .in1(N__1875),
            .in2(_gnd_net_),
            .in3(N__1869),
            .lcout(rst_cntZ0Z_5),
            .ltout(),
            .carryin(un1_rst_cnt_1_cry_4),
            .carryout(un1_rst_cnt_1_cry_5),
            .clk(N__2370),
            .ce(),
            .sr(N__1982));
    defparam rst_cnt_6_LC_2_7_6.C_ON=1'b1;
    defparam rst_cnt_6_LC_2_7_6.SEQ_MODE=4'b1000;
    defparam rst_cnt_6_LC_2_7_6.LUT_INIT=16'b0110011011001100;
    LogicCell40 rst_cnt_6_LC_2_7_6 (
            .in0(N__2331),
            .in1(N__1866),
            .in2(_gnd_net_),
            .in3(N__1860),
            .lcout(rst_cntZ0Z_6),
            .ltout(),
            .carryin(un1_rst_cnt_1_cry_5),
            .carryout(un1_rst_cnt_1_cry_6),
            .clk(N__2370),
            .ce(),
            .sr(N__1982));
    defparam rst_cnt_7_LC_2_7_7.C_ON=1'b1;
    defparam rst_cnt_7_LC_2_7_7.SEQ_MODE=4'b1000;
    defparam rst_cnt_7_LC_2_7_7.LUT_INIT=16'b0110011011001100;
    LogicCell40 rst_cnt_7_LC_2_7_7 (
            .in0(N__2324),
            .in1(N__1857),
            .in2(_gnd_net_),
            .in3(N__1851),
            .lcout(rst_cntZ0Z_7),
            .ltout(),
            .carryin(un1_rst_cnt_1_cry_6),
            .carryout(un1_rst_cnt_1_cry_7),
            .clk(N__2370),
            .ce(),
            .sr(N__1982));
    defparam rst_cnt_8_LC_2_8_0.C_ON=1'b1;
    defparam rst_cnt_8_LC_2_8_0.SEQ_MODE=4'b1000;
    defparam rst_cnt_8_LC_2_8_0.LUT_INIT=16'b0110011011001100;
    LogicCell40 rst_cnt_8_LC_2_8_0 (
            .in0(N__2327),
            .in1(N__1848),
            .in2(_gnd_net_),
            .in3(N__1842),
            .lcout(rst_cntZ0Z_8),
            .ltout(),
            .carryin(bfn_2_8_0_),
            .carryout(un1_rst_cnt_1_cry_8),
            .clk(N__2368),
            .ce(),
            .sr(N__1981));
    defparam rst_cnt_9_LC_2_8_1.C_ON=1'b1;
    defparam rst_cnt_9_LC_2_8_1.SEQ_MODE=4'b1000;
    defparam rst_cnt_9_LC_2_8_1.LUT_INIT=16'b0110011011001100;
    LogicCell40 rst_cnt_9_LC_2_8_1 (
            .in0(N__2320),
            .in1(N__1839),
            .in2(_gnd_net_),
            .in3(N__1833),
            .lcout(rst_cntZ0Z_9),
            .ltout(),
            .carryin(un1_rst_cnt_1_cry_8),
            .carryout(un1_rst_cnt_1_cry_9),
            .clk(N__2368),
            .ce(),
            .sr(N__1981));
    defparam rst_cnt_10_LC_2_8_2.C_ON=1'b1;
    defparam rst_cnt_10_LC_2_8_2.SEQ_MODE=4'b1000;
    defparam rst_cnt_10_LC_2_8_2.LUT_INIT=16'b0110011011001100;
    LogicCell40 rst_cnt_10_LC_2_8_2 (
            .in0(N__2325),
            .in1(N__1830),
            .in2(_gnd_net_),
            .in3(N__1824),
            .lcout(rst_cntZ0Z_10),
            .ltout(),
            .carryin(un1_rst_cnt_1_cry_9),
            .carryout(un1_rst_cnt_1_cry_10),
            .clk(N__2368),
            .ce(),
            .sr(N__1981));
    defparam rst_cnt_11_LC_2_8_3.C_ON=1'b1;
    defparam rst_cnt_11_LC_2_8_3.SEQ_MODE=4'b1000;
    defparam rst_cnt_11_LC_2_8_3.LUT_INIT=16'b0110011011001100;
    LogicCell40 rst_cnt_11_LC_2_8_3 (
            .in0(N__2318),
            .in1(N__1821),
            .in2(_gnd_net_),
            .in3(N__1815),
            .lcout(rst_cntZ0Z_11),
            .ltout(),
            .carryin(un1_rst_cnt_1_cry_10),
            .carryout(un1_rst_cnt_1_cry_11),
            .clk(N__2368),
            .ce(),
            .sr(N__1981));
    defparam rst_cnt_12_LC_2_8_4.C_ON=1'b1;
    defparam rst_cnt_12_LC_2_8_4.SEQ_MODE=4'b1000;
    defparam rst_cnt_12_LC_2_8_4.LUT_INIT=16'b0110011011001100;
    LogicCell40 rst_cnt_12_LC_2_8_4 (
            .in0(N__2326),
            .in1(N__1812),
            .in2(_gnd_net_),
            .in3(N__1806),
            .lcout(rst_cntZ0Z_12),
            .ltout(),
            .carryin(un1_rst_cnt_1_cry_11),
            .carryout(un1_rst_cnt_1_cry_12),
            .clk(N__2368),
            .ce(),
            .sr(N__1981));
    defparam rst_cnt_13_LC_2_8_5.C_ON=1'b1;
    defparam rst_cnt_13_LC_2_8_5.SEQ_MODE=4'b1000;
    defparam rst_cnt_13_LC_2_8_5.LUT_INIT=16'b0110011011001100;
    LogicCell40 rst_cnt_13_LC_2_8_5 (
            .in0(N__2319),
            .in1(N__2034),
            .in2(_gnd_net_),
            .in3(N__2028),
            .lcout(rst_cntZ0Z_13),
            .ltout(),
            .carryin(un1_rst_cnt_1_cry_12),
            .carryout(un1_rst_cnt_1_cry_13),
            .clk(N__2368),
            .ce(),
            .sr(N__1981));
    defparam un1_rst_cnt_1_cry_13_c_THRU_CRY_0_LC_2_8_6.C_ON=1'b1;
    defparam un1_rst_cnt_1_cry_13_c_THRU_CRY_0_LC_2_8_6.SEQ_MODE=4'b0000;
    defparam un1_rst_cnt_1_cry_13_c_THRU_CRY_0_LC_2_8_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_rst_cnt_1_cry_13_c_THRU_CRY_0_LC_2_8_6 (
            .in0(_gnd_net_),
            .in1(N__2024),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_rst_cnt_1_cry_13),
            .carryout(un1_rst_cnt_1_cry_13_THRU_CRY_0_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam un1_rst_cnt_1_cry_13_c_THRU_CRY_1_LC_2_8_7.C_ON=1'b1;
    defparam un1_rst_cnt_1_cry_13_c_THRU_CRY_1_LC_2_8_7.SEQ_MODE=4'b0000;
    defparam un1_rst_cnt_1_cry_13_c_THRU_CRY_1_LC_2_8_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 un1_rst_cnt_1_cry_13_c_THRU_CRY_1_LC_2_8_7 (
            .in0(_gnd_net_),
            .in1(N__2025),
            .in2(GNDG0),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(un1_rst_cnt_1_cry_13_THRU_CRY_0_THRU_CO),
            .carryout(un1_rst_cnt_1_cry_13_THRU_CRY_1_THRU_CO),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam rst_cnt_esr_14_LC_2_9_0.C_ON=1'b0;
    defparam rst_cnt_esr_14_LC_2_9_0.SEQ_MODE=4'b1000;
    defparam rst_cnt_esr_14_LC_2_9_0.LUT_INIT=16'b0011001111001100;
    LogicCell40 rst_cnt_esr_14_LC_2_9_0 (
            .in0(_gnd_net_),
            .in1(N__2010),
            .in2(_gnd_net_),
            .in3(N__2013),
            .lcout(rst_cntZ0Z_14),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2371),
            .ce(N__1995),
            .sr(N__1983));
    defparam LED2_obuf_RNO_LC_4_2_3.C_ON=1'b0;
    defparam LED2_obuf_RNO_LC_4_2_3.SEQ_MODE=4'b0000;
    defparam LED2_obuf_RNO_LC_4_2_3.LUT_INIT=16'b1011101110001000;
    LogicCell40 LED2_obuf_RNO_LC_4_2_3 (
            .in0(N__2175),
            .in1(N__1929),
            .in2(_gnd_net_),
            .in3(N__1959),
            .lcout(LED2_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam LED1_obuf_RNO_LC_4_2_4.C_ON=1'b0;
    defparam LED1_obuf_RNO_LC_4_2_4.SEQ_MODE=4'b0000;
    defparam LED1_obuf_RNO_LC_4_2_4.LUT_INIT=16'b1101110110001000;
    LogicCell40 LED1_obuf_RNO_LC_4_2_4 (
            .in0(N__1928),
            .in1(N__2181),
            .in2(_gnd_net_),
            .in3(N__1905),
            .lcout(LED1_c),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_1_LC_4_6_0.C_ON=1'b0;
    defparam clk_div_1_LC_4_6_0.SEQ_MODE=4'b1000;
    defparam clk_div_1_LC_4_6_0.LUT_INIT=16'b1010010101011010;
    LogicCell40 clk_div_1_LC_4_6_0 (
            .in0(N__2113),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2133),
            .lcout(clk_divZ0Z_1),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2378),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_0_LC_4_6_1.C_ON=1'b0;
    defparam clk_div_0_LC_4_6_1.SEQ_MODE=4'b1000;
    defparam clk_div_0_LC_4_6_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 clk_div_0_LC_4_6_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2112),
            .lcout(clk_divZ0Z_0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2378),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNI91U1_1_LC_4_7_0.C_ON=1'b1;
    defparam clk_div_RNI91U1_1_LC_4_7_0.SEQ_MODE=4'b0000;
    defparam clk_div_RNI91U1_1_LC_4_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNI91U1_1_LC_4_7_0 (
            .in0(_gnd_net_),
            .in1(N__2131),
            .in2(N__2114),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_7_0_),
            .carryout(clk_div_2_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNIF3T2_2_LC_4_7_1.C_ON=1'b1;
    defparam clk_div_RNIF3T2_2_LC_4_7_1.SEQ_MODE=4'b0000;
    defparam clk_div_RNIF3T2_2_LC_4_7_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNIF3T2_2_LC_4_7_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2088),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_1),
            .carryout(clk_div_2_cry_2),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNIM6S3_3_LC_4_7_2.C_ON=1'b1;
    defparam clk_div_RNIM6S3_3_LC_4_7_2.SEQ_MODE=4'b0000;
    defparam clk_div_RNIM6S3_3_LC_4_7_2.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNIM6S3_3_LC_4_7_2 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2070),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_2),
            .carryout(clk_div_2_cry_3),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNIUAR4_4_LC_4_7_3.C_ON=1'b1;
    defparam clk_div_RNIUAR4_4_LC_4_7_3.SEQ_MODE=4'b0000;
    defparam clk_div_RNIUAR4_4_LC_4_7_3.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNIUAR4_4_LC_4_7_3 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2052),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_3),
            .carryout(clk_div_2_cry_4),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNI7GQ5_5_LC_4_7_4.C_ON=1'b1;
    defparam clk_div_RNI7GQ5_5_LC_4_7_4.SEQ_MODE=4'b0000;
    defparam clk_div_RNI7GQ5_5_LC_4_7_4.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNI7GQ5_5_LC_4_7_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2520),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_4),
            .carryout(clk_div_2_cry_5),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNIHMP6_6_LC_4_7_5.C_ON=1'b1;
    defparam clk_div_RNIHMP6_6_LC_4_7_5.SEQ_MODE=4'b0000;
    defparam clk_div_RNIHMP6_6_LC_4_7_5.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNIHMP6_6_LC_4_7_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2502),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_5),
            .carryout(clk_div_2_cry_6),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNISTO7_7_LC_4_7_6.C_ON=1'b1;
    defparam clk_div_RNISTO7_7_LC_4_7_6.SEQ_MODE=4'b0000;
    defparam clk_div_RNISTO7_7_LC_4_7_6.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNISTO7_7_LC_4_7_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2484),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_6),
            .carryout(clk_div_2_cry_7),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNI86O8_8_LC_4_7_7.C_ON=1'b1;
    defparam clk_div_RNI86O8_8_LC_4_7_7.SEQ_MODE=4'b0000;
    defparam clk_div_RNI86O8_8_LC_4_7_7.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNI86O8_8_LC_4_7_7 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2466),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_7),
            .carryout(clk_div_2_cry_8),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNILFN9_9_LC_4_8_0.C_ON=1'b1;
    defparam clk_div_RNILFN9_9_LC_4_8_0.SEQ_MODE=4'b0000;
    defparam clk_div_RNILFN9_9_LC_4_8_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNILFN9_9_LC_4_8_0 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(N__2448),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_4_8_0_),
            .carryout(clk_div_2_cry_9),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNIAAMP_10_LC_4_8_1.C_ON=1'b1;
    defparam clk_div_RNIAAMP_10_LC_4_8_1.SEQ_MODE=4'b0000;
    defparam clk_div_RNIAAMP_10_LC_4_8_1.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_RNIAAMP_10_LC_4_8_1 (
            .in0(_gnd_net_),
            .in1(N__2426),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(clk_div_2_cry_9),
            .carryout(clk_div_2_cry_10),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_RNI06L91_11_LC_4_8_2.C_ON=1'b0;
    defparam clk_div_RNI06L91_11_LC_4_8_2.SEQ_MODE=4'b0000;
    defparam clk_div_RNI06L91_11_LC_4_8_2.LUT_INIT=16'b0011001111001100;
    LogicCell40 clk_div_RNI06L91_11_LC_4_8_2 (
            .in0(_gnd_net_),
            .in1(N__2192),
            .in2(_gnd_net_),
            .in3(N__2217),
            .lcout(clk_div_RNI06L91Z0Z_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_11_LC_4_8_5.C_ON=1'b0;
    defparam clk_div_11_LC_4_8_5.SEQ_MODE=4'b1000;
    defparam clk_div_11_LC_4_8_5.LUT_INIT=16'b1111111100000000;
    LogicCell40 clk_div_11_LC_4_8_5 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2210),
            .lcout(clk_div_i_11),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2372),
            .ce(),
            .sr(_gnd_net_));
    defparam LED1_m0_r_LC_5_2_1.C_ON=1'b0;
    defparam LED1_m0_r_LC_5_2_1.SEQ_MODE=4'b1000;
    defparam LED1_m0_r_LC_5_2_1.LUT_INIT=16'b0000000011111111;
    LogicCell40 LED1_m0_r_LC_5_2_1 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2396),
            .lcout(LED1_m0_rZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2381),
            .ce(N__2270),
            .sr(_gnd_net_));
    defparam LED2_m0_r_LC_5_2_4.C_ON=1'b0;
    defparam LED2_m0_r_LC_5_2_4.SEQ_MODE=4'b1000;
    defparam LED2_m0_r_LC_5_2_4.LUT_INIT=16'b0000000011111111;
    LogicCell40 LED2_m0_r_LC_5_2_4 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2147),
            .lcout(LED2_m0_rZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2381),
            .ce(N__2270),
            .sr(_gnd_net_));
    defparam BUT2_r_LC_5_2_6.C_ON=1'b0;
    defparam BUT2_r_LC_5_2_6.SEQ_MODE=4'b1000;
    defparam BUT2_r_LC_5_2_6.LUT_INIT=16'b1111111100000000;
    LogicCell40 BUT2_r_LC_5_2_6 (
            .in0(_gnd_net_),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(N__2169),
            .lcout(BUT2_rZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2381),
            .ce(N__2270),
            .sr(_gnd_net_));
    defparam clk_div_1_cry_1_c_LC_5_7_0.C_ON=1'b1;
    defparam clk_div_1_cry_1_c_LC_5_7_0.SEQ_MODE=4'b0000;
    defparam clk_div_1_cry_1_c_LC_5_7_0.LUT_INIT=16'b0000000000000000;
    LogicCell40 clk_div_1_cry_1_c_LC_5_7_0 (
            .in0(_gnd_net_),
            .in1(N__2132),
            .in2(N__2115),
            .in3(_gnd_net_),
            .lcout(),
            .ltout(),
            .carryin(bfn_5_7_0_),
            .carryout(clk_div_1_cry_1),
            .clk(_gnd_net_),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_2_LC_5_7_1.C_ON=1'b1;
    defparam clk_div_2_LC_5_7_1.SEQ_MODE=4'b1000;
    defparam clk_div_2_LC_5_7_1.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_2_LC_5_7_1 (
            .in0(_gnd_net_),
            .in1(N__2087),
            .in2(_gnd_net_),
            .in3(N__2073),
            .lcout(clk_divZ0Z_2),
            .ltout(),
            .carryin(clk_div_1_cry_1),
            .carryout(clk_div_1_cry_2),
            .clk(N__2379),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_3_LC_5_7_2.C_ON=1'b1;
    defparam clk_div_3_LC_5_7_2.SEQ_MODE=4'b1000;
    defparam clk_div_3_LC_5_7_2.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_3_LC_5_7_2 (
            .in0(_gnd_net_),
            .in1(N__2069),
            .in2(_gnd_net_),
            .in3(N__2055),
            .lcout(clk_divZ0Z_3),
            .ltout(),
            .carryin(clk_div_1_cry_2),
            .carryout(clk_div_1_cry_3),
            .clk(N__2379),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_4_LC_5_7_3.C_ON=1'b1;
    defparam clk_div_4_LC_5_7_3.SEQ_MODE=4'b1000;
    defparam clk_div_4_LC_5_7_3.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_4_LC_5_7_3 (
            .in0(_gnd_net_),
            .in1(N__2051),
            .in2(_gnd_net_),
            .in3(N__2037),
            .lcout(clk_divZ0Z_4),
            .ltout(),
            .carryin(clk_div_1_cry_3),
            .carryout(clk_div_1_cry_4),
            .clk(N__2379),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_5_LC_5_7_4.C_ON=1'b1;
    defparam clk_div_5_LC_5_7_4.SEQ_MODE=4'b1000;
    defparam clk_div_5_LC_5_7_4.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_5_LC_5_7_4 (
            .in0(_gnd_net_),
            .in1(N__2519),
            .in2(_gnd_net_),
            .in3(N__2505),
            .lcout(clk_divZ0Z_5),
            .ltout(),
            .carryin(clk_div_1_cry_4),
            .carryout(clk_div_1_cry_5),
            .clk(N__2379),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_6_LC_5_7_5.C_ON=1'b1;
    defparam clk_div_6_LC_5_7_5.SEQ_MODE=4'b1000;
    defparam clk_div_6_LC_5_7_5.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_6_LC_5_7_5 (
            .in0(_gnd_net_),
            .in1(N__2501),
            .in2(_gnd_net_),
            .in3(N__2487),
            .lcout(clk_divZ0Z_6),
            .ltout(),
            .carryin(clk_div_1_cry_5),
            .carryout(clk_div_1_cry_6),
            .clk(N__2379),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_7_LC_5_7_6.C_ON=1'b1;
    defparam clk_div_7_LC_5_7_6.SEQ_MODE=4'b1000;
    defparam clk_div_7_LC_5_7_6.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_7_LC_5_7_6 (
            .in0(_gnd_net_),
            .in1(N__2483),
            .in2(_gnd_net_),
            .in3(N__2469),
            .lcout(clk_divZ0Z_7),
            .ltout(),
            .carryin(clk_div_1_cry_6),
            .carryout(clk_div_1_cry_7),
            .clk(N__2379),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_8_LC_5_7_7.C_ON=1'b1;
    defparam clk_div_8_LC_5_7_7.SEQ_MODE=4'b1000;
    defparam clk_div_8_LC_5_7_7.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_8_LC_5_7_7 (
            .in0(_gnd_net_),
            .in1(N__2465),
            .in2(_gnd_net_),
            .in3(N__2451),
            .lcout(clk_divZ0Z_8),
            .ltout(),
            .carryin(clk_div_1_cry_7),
            .carryout(clk_div_1_cry_8),
            .clk(N__2379),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_9_LC_5_8_0.C_ON=1'b1;
    defparam clk_div_9_LC_5_8_0.SEQ_MODE=4'b1000;
    defparam clk_div_9_LC_5_8_0.LUT_INIT=16'b1001100101100110;
    LogicCell40 clk_div_9_LC_5_8_0 (
            .in0(_gnd_net_),
            .in1(N__2447),
            .in2(_gnd_net_),
            .in3(N__2433),
            .lcout(clk_divZ0Z_9),
            .ltout(),
            .carryin(bfn_5_8_0_),
            .carryout(clk_div_1_cry_9),
            .clk(N__2374),
            .ce(),
            .sr(_gnd_net_));
    defparam clk_div_10_LC_5_8_1.C_ON=1'b0;
    defparam clk_div_10_LC_5_8_1.SEQ_MODE=4'b1000;
    defparam clk_div_10_LC_5_8_1.LUT_INIT=16'b0011001111001100;
    LogicCell40 clk_div_10_LC_5_8_1 (
            .in0(_gnd_net_),
            .in1(N__2427),
            .in2(_gnd_net_),
            .in3(N__2430),
            .lcout(clk_divZ0Z_10),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2374),
            .ce(),
            .sr(_gnd_net_));
    defparam BUT1_r_LC_6_2_2.C_ON=1'b0;
    defparam BUT1_r_LC_6_2_2.SEQ_MODE=4'b1000;
    defparam BUT1_r_LC_6_2_2.LUT_INIT=16'b1010101010101010;
    LogicCell40 BUT1_r_LC_6_2_2 (
            .in0(N__2415),
            .in1(_gnd_net_),
            .in2(_gnd_net_),
            .in3(_gnd_net_),
            .lcout(BUT1_rZ0),
            .ltout(),
            .carryin(_gnd_net_),
            .carryout(),
            .clk(N__2382),
            .ce(N__2271),
            .sr(_gnd_net_));
endmodule // led_but_ex1
